PK   �K�XЪ^-�&  kv    cirkitFile.json�[��Hr�JC~9(�3��K������6v��Cw��x���j��R�ō��ΠT7^$����a���t��׏�`0#��u�/n�E��7����~�ۮn(�Z}.��/�˿5W��Ͷ8슿�˻ϫ�������]��MY�w�M�*Ɍ�����ȥq�&+��J�j�m�ia
�������
$V0��
���RSX1�T�N� U0E"f�*�"3HL���
���RSx1�T!�(y�K
@���J�K�D���K�D��L�D���L�D��M�D���M�D��N�D���N�D�[q�{�����}���/P��n����[�m��v��q8��a�D� tZ�W����Tt7�E�øX"P�øX"P�øX"P�øX"P�øX"P��ЕCC����_	b���ʻ��HC��.+�%��- ���y��0.��0.��0t�����`��D����m.]V��o��)��- ��0.��0.�0�Xb
+t��t/0��a�!��%�wb�Thʐ�
/B��K
�{C,(�_,a�D���B���B���B���B���0)��<�%�<v�%�t&y1s���2�<'�8,�0E*�O�#�<����I<T�/w�m�=~��mT�k�u�E��M���js��օ�ߗ�_i,����,w	��I{}1"9v0�a�Kg� �v�����t�����������k;�����t!����am�#,]�am�`m�#,]�(`m�bm�#,�)2��2��t��3E��]�����t��X�y��t���/p��cpf��#0;�:�@�����	�3,���{m���Y���|��9�~�L�G`>�Fl?p���#0��8������%���:�|��`��3,��x-�~���G`�׋P ̃��d�(6�i_�\��\��%�/X>��b!���$�p��ӗ��`���+����/X>���0�������|��l?p���#0�����`���z! �~��@�}̥�Gp�3�<����O�~�|����OD��/X>��ZQ�������|��l?p���#0������#/p�b���/X>��h�������|�cC�7H$�G�
���ˣ�����Xp���#0/��<y��#0�����`��Ǖ��s���G`>�� �8}�����;��N_�|��`���,���$�~�e*�u*��Ł�N_�|��:"`��g_�|��&`���,����
�~���G`>.�8������`헀�,���TO��Yma}+�o��S���� ��.	8u����++�\����z���Ӄ���$��G`>.��z�>z�>8�I�YO�z�|���c`���,���U�d�|����8�&,�x�� )ysO�	�k��F#�&3U
η�u�dOR*]���<�<����E)8������ ��ι�|t��9�%y�����Q��F�N�]���Yf�x�!��������7.lޯ���y������������.lޯ��y�(����j�K�F�vB�쨸�����.m/���΁K��o�[���B��j���4�	�o�����B�l��������-m/����^K_\B�섵����+����QK��o�����B�l������-m/����;���vII_O,�Y����P�v��+!ؕ8)JoPD�2\f5��-3K�};�������V6�}����,������j��J��䃳�OǅYͧ�yV�鷒u�ViKQ��8rM�F�Y�4�^���̵�j>}�O_���g�����$��:k"�l������6�|bJ���9��\���g�}N������]Q�nw���Wɨc���L���J�8���C2|�0D !Î�!	~�a�@B��n"���&�$d��!	����b�@B�U�H\�ƅmX�&X�F)�nD����(%Ӎ���`�`�d�j,�,���L7�b��񸋾��?|�KX�aq�d�YS�Ԇ$[���(%��v��`q<��q���fe@L�8��8J�����O�8��8J�t�\�t��F _���	�QJ���1�FRpC)�8naq�d��H,���,,�[XG)�n�tRJ�y+d��q���f�A�������q���f�AL�8�`q�QI��7(�P���(%�� cJQ����q���1����QJ�6���	,���x�5�	�XG)�
_nv7�	��	,���xu'�	Ǔ.����	�XG)u+�@�]
��),��\[��`q���c�WL�?S�E��v+����J*���Q����J*���]����J*��������J*�!�R�k�T�����A*v헐�X@��TXCEŮ��2h��
�)��f�@�j��
�)�Ud�@�j��
�)�%b�@�j��
+���d\*��C��6��V)�RJ�t�.�I�H'�R�%Z��\Ƕ:ٗ
-���7�:����ThI����ױ�N�BK:���AǶ:��
-���Z��dc*��C�kJtl����В-��ѱ�NV�BK:���Ggba���I�0�����B�����:y�
-���+�*͈)M���e�N^��e*��C�k�tl����В-��ӱ�N^�BK:��&QǶ:y�
-����J���e*��C�kDul;�t �[��l�b��,���ThI�����|��3_�BK:���XǶ:y�
-���j���e*��C�k�ul������:y���ˬN^�BK:��6_Ƕ:y�
-��r��3D�V���h!F��ˬN^�BK:�\�AǶ:�e*��C˵+tl����В-��P�����ThI��k���V'/S�%Z���c[��L��th����mu�2Zҡ�5:�UZI���L'/s:y����ThI��k��Vg�L��th����mu�2Zҡ�N:����ThI��kQ��V'/S�%Z���b�D'/S�%���r7cŁd�H���e*�\�L�ou�2Zҡ���[��l�-���N^���e*��C˵�tl�T�C�̇N^���e�N^�BK:�\�PǶ:y�
-��rMF�w�N^6B��E�V'/���CW��1Z�R��,�Y_�BKc�#�̗�:y�
-��r�R���e*�4��y��$oҼ]�Q;�\U���i��45>�lO�üPe���B����U&�x/T����Pe�V�B����U&�Q/T�� �Pe���R�9/�{�6}]*��ߩ�U��`<xjӥ2��&t�Ƌ�6�\*��/�ڥr�Ƌ���\*�����`�xj_åo]�O��Tԕ�x�ԶzKe0^<�y�R�Om6�T��S�-��x��vg�2~��mT�k�u�E��M���js����.�p㈅*4>ƵPsE��Ƈ)�\|(g�\|&g�t��p;�g���B��F��C���+������j��J�/���T.>�T.��,��a�:j�����y��n#�MS��m}s�.�T.�e��E��R�l
�͓�ꬉ��U�c�:��$�)]<�.sT.�e��e��Qyi��;��+��Y�|}�]���j�<���K��[LgwH�t�B2�?@�@B�{wA�@B�{B�@B�{�B�@B�{?C�@B�΃��L74!	��0#&D�6.l��6�7J�GS1L��M���R2�q^,~,����q����(%s�0��x��(%s��0��߸8,�ǰ8�R2��	,�ǰ8�R2�i,�ǰ8�R2�	,�ǰ8�R2ǩ&L:���QJ�8	�a���R`q���8J���0L�8naq�d���&X��8�R2��Q,�;XG)���-�	�,����
�	7&���q��(%.Zc��q��(%.� c��q��(%^�������QJ����	,���x�1�	7���ބ���QJ�8���	,���x1"�	�SXG)��7,���8>��|!�`�$Z����J*���j��"I�*Ю���j��I�*Ю���j�A��*Ю����.���@,��J*���b�A��4XI�5�QT�:�S��+���bP��
��+���bP��
��+���bP��
��+���7�:��NƥBK:��m��m��.��K'�"�ċt2/Zҡ�o�ul��}�В-3�c[�L��th����da*��C�ktl����В-��б�N6�BK:���DǶ:�
-������de*��C�k|t&t�2Zҡ�J:����ThI���\��ViFLiJL'/�u�X'/S�%Z^�c[��L��thy-��mu�2Zҡ�5�:����ThI���V��V'/S�%Z^#�c[��L��thy���mu�2Zҡ�5�:&��e*��C�k�ul����В-��ֱ�N^�BK:��\ǶJ_+*}����Y�����e*��C�k�ul����В-�б�N^�BK:�\+AǶ:y�
-��r����e*��C˵+tl����В-��P�����ThI��k���V'/S�%Z���c[��L��th����mu�2Zҡ�5:�UZI���L'/s:y����ThI��k��V'/S�%Z�}�c[��L��th����mu�2Zҡ�ZT:����ThI��kj��6���ThI��k���V'/S�%Z�q�c[��L��th�V��mu�2Zҡ�s:����ThI��k���V�ʇR���,�����L��th����mu�2Zҡ嚌:����ThI��kK��V'/S�%Z���b�T'/S�%Z���c[��L��th�f��mu�2Z�G��Ut�7iޮ�(�E��m�봎�u��e6�'�a^�2Q�v��D5م*u��LT�^�2Q+{��Du�*���LT�^�2Q�y�ׁ��S��.�����֪Ke0<���R�Om�T��S�q.��`�O�R�T��S{A.��x�Ԏ�Ke0^<���ҷ.Ƌ�v\*�J`�xj[��2/�ڼn�Ƌ���[*��⩍ؖ�`�xj��g�vY��6*׵�ܺ΢��&J|S����k��]�Y*/i�
�.>��T.>��T.>��T.>��T.>�m��敍b��D3nW_GUI�f��_��Y*�e��E��r�_���J[�Z�Ǒk�6�ޘ�ڤ1����7��2K�]f�\��,��v�`�<	q�Κ�9[E>�>��M2����3�2G�]�\����v��*�篇�����Ŧ�uu�^�~�������l�ݾn�����MI�٧+ѯ'9vJ���kɛK�B(+�IݎK�׃��I����/�M�K	��@n�TF�{���_{'�1�[���1R�~e9N�fI�(�y=i �Mj~÷�Me��q��o���G�7�
��>=v��͗�ϡ�Tn��Ӈ N�ǿ���o��oڇ�@���#T߸G�!Bv�wN޿�@������ `� i�� r�cOa0T�LBOh:�o��Uy��+�;�c�o�vE����ݓQ	o]�Y�Pű0�'���O�!T�CO��* <l����P���ӟwm{���+6�����r
�[Z,a�� !�X�tSIB
��馢�b	�M�)���jR�%L7U/�K�n�_H!�0���B
���&R�%��kdi�BDOD��OP��9~P-� �PQ��9~�-� �QR��9~T.� �RS��9~�.� ���x��"V�1 ��5��C})G<0�ɅX�h+�0ǕR@���V�a�k��h��\�WO���b�o�rs\�!�;��dB,@�k���)bt 1< ��m��DF�������{! �Z@�k��)�0���9."�b��_��9.c�r ��D[�W pX��:�謃�� �5�F3�c$�%��r.� �| ��5��,`�|@�kp�R  �&��+���� �db6^@x�kpYB  �&#�R�e�	 ��5��������h��m�ѻ�D���� �OB��2(�W��u�Dz�#0�)��pz�a��g�Ay=��~X>�bP������|!W�oP�\x�X>���~��������/t���^/���|����A��#0�)��qz�a��g�A�p��~X>���4:��?E�����tB�D�Й��Є�y.چ�lLHhB��mCtF&$4!��!:+��?�F����		Mȟ��m��N���&�O��6Dg(`BB�2 ��Y
��Є���b�Y@o��d ����%F�-`BB�@16�Ϡ�Ӗ����LHhB^���!:m����m�N[���&�Qh��0!�	y]چ�LHh��i06$�V��iXjt��0!�	�Ů����E�i��.�m�N[���&�E�h��0!�	y�(چ�o�����N[,:m���m�N[���&|]Uc�AR��l�-��b��R����b���&Vl�
bl�N[���mCt�&$4!���С�0!�	� چ�LHhB�^��!:m��+/�m�N[���&�2h��׭���N[:m���q�m��m�����m��S���&��'h��0!�	�hچ�<LHhB.8�a��S���&n�6��8}�I�i���������		M8��p���t3
bL��bt&$4!��B�� ���$�,&Ag1`BBr�.��Y��Єíz����cL�Nj���wPĸ� e��"Q7���4,�@��q�{g��)��``�Z =5��s0!�	��چ�LH����M�&��u%���U��|��Q�NS�̦��f���..l?(���������:���.l?�����������¤�
�.��J=p�C�R���[* ���.lK�~8��l����[�-�B�'��Z* ���FWK��8�Zj�����7-}�I=q�A�R�kY�ý��
H=q�]�R�'7�Y* ���4K��8���Y��]�����um"���(w���Tm�}�ں�V��F*��9���e�{Ȑ���<��ڟyg�φ�q�rm���F��C�_,������j��J���J�ڟyf�?�,�ڟ���Q[�-E����5uyoLdmҘzml�s�?���������j��)�/OB�&r�V�����<o��'�t��������i���?^��W��v��8� x������W7V<4ǣ�8��C�A����=�xc%^iҭN�*�ta��\Ⓣ�&>��|��-bnw��"�1���E�-bns��[Xna���p����[Xna����[8n�Ex�|
�3B��Bs¡�'���g������w~���� 7�xM���M�@gF���+B����_0��R:B��:'��ݮ$�7�(�� Ȍ �B ��+��2�P��	��,�K�D(v#'C(#_�hj8�5 $q����I:�C�y��l*�_m��~�;_P�b'CB�+4�`�zߋW����Pܖ��{ �{�]��h�8��ŧC��=��C�t�%�C��Pz:�e�C��P~:���!38D��E#�O���٣"�H>Y���]��/<`�mw�����.2�v������?4E�����?��m��������+O!��_�C��v�~��k��Mӥ_��/v�`���~��8�-���������������w���vxW��?�~���� ��i���&�o���oַ�����~���M?�`�/���-��þٟ����=�����[7��o��o 8�'t�6��.�����(N��Fͮr�]'&3�����?�U�Vyc�:jېTx��Qkc�T�M�$6�R����f��]�BZw(��QhVrw���7A�<®n����}uۜn�p�ur���W�ꧫ6�+�6s�k����||<-�6;͙��?ɍ�����,;~�=��gŒ�X<~8�^�O\��O*'+�I�ǻk��?�x7~<�c��0�����l��;6��	r�����Ξ��l���D���������΢���b�"��Y�ʋ�K^O^�J|���QG�w쬗V=�d{w��=<��ѳ�]i�0�!y�ϣǟ��ý�*s�=>�t���|�:��1~V/ MܯA8?���J�g�rv�G眝�Ι�y~jo��ݧ��^�0I�U������׏�K�������o͡��qu�q����I��iŶl#W�,�1E.ueK�pҝ��zw�o�;|���ض1��U�D��$r�������)���׭�|ז�E��ʓ�I�(d1u�ț(�3WW�K��ϟ����{8�hL�l]�m���e�Zz�#JJ�M�Y�6���q��%�l����|%����/���-�YRF��Y�b�2N��MU�d���+S|_���ß���8k�����ok����&��u<)�U���|��o^�G���T���	]���J:u��5��q���u��w�n�w[�߅��f���{�?��z�)����˺�o�6ծk����x���G����?�����?����\�\���fĽ�C�W.�J���SIR��n�˫4�K۬�:�K�\,�*M"�.X���O�VQp�uޖ�^�d�����-��.�ΦvQ�[��	�gS�U��t1���m誅.f��:�>�F�M�8t��v��w���Ǐ��w���}sx��?���׏�����?�?�����x����s�o��v���w����	g������N�v���Rn�#2��)M}��K�#�O�mS:���2W�c��w�-�Ow|���uȠ(;�|�O]W�o��O��z�{�ˮ��^��1#)���uP��B��O���*I�k:���E�_��}R�2�&��v�;ʪ�$��:	�G�r�w�z׳&f�����U���5t�P����P�x 6׉�yb����ػ��%z����5����F��N{�Kc���;8�-wuQ������s݀ݷ��+���a�C$�OO�0N�|�g/�g��!.�Y��s���4
Al�$k�eUm�Y����O?�<:�����<K�#��}�C��o�>��Gϊ�Mn�K_e)�~�އ�<�������~ݬ�j�u\GY钨��:j,eq^�T�Y�7kRt���n����H߯�#�%�;�u���x��|��}�����t>:��&I�i�@Ҽ]<�GyZ֞Lȉ�z��͙X��|�q�,����q��_��O���F���p��a[w�u؅��r�}$�}�uA����:���eS>�{$��6w�4����Q��:�Ҕ��5��6gRV����������p��/���
������r/7t׻n�?��_X׵7cx�ٞ:Ӣ��i�����i��_~���?����~���U�n��ޗ�ϝx�
>�x��O�{>�S������|��=�<�S��e���F�ʒ�w֧�C�f�,�0{���&V���]x�_�	E�����Y��St�ON1�o�:�:��:�:#�K]�17��9��5�ǁ�K��;k���Ƙ���v���3��s)��L���）u�����n�O�7����e��J�����;�ql#;�P�-��;ԹW������e��P�,W靕�:����^n�[�D�q���:o�ng�u���Q�������]�ٓ�BG��9�-���o8���}���;�no�{��F�.���Y�q �o9k��m���m��<����{>�I��<~V?���)�-g͍<���w<R���<���Fj��S�1��} ?g��wV���k�p��ߠc�m��濉�n��.��u�ʱki��g��x��p��1v��>��z�#��A;���nk�:v��ˣw�7u�;��[ۡ� ��0����q��Y��������{?�w y���9���xrs{������o�[.�|������������n���C�?�����n��Mu����o�N����PK   J�X�R�� $� /   images/179c08ce-6e18-4019-8002-932a24469ad1.png�z�[�a�>XJ(*�"���� A�P:��0�]"�HHwwMb��Cr��l�6`�o�}�?�w]_.v}ೋ�9�<�}��|X�k-eJ

JU��:$$��HHn�ݼA�S����p�榠�w���w���wrgc7�⋴�NO�p��������{w���	�s�YY:�8�ڦ�dHH���|�畱��s7���8Yp+��~b��x#�񋈻�jIPH�i43l�q�Ͳ�SĚ�4"^6^DRd+>�[��:�[�WJ���=I�)�C+Ocy�;?(���(�x��ZBD�$��#�e�0,Y�[曽�t?'��|ߌ�D��Y��2���I�o͕7`�6`�Ü	�����`���C(�͚ɀS�@��2�͸�H���j�~2��g��s������n���������:�#���9rHC4�NM]O�~Kˌ�S8_>��C���d�K%I�:���*E�J�<��:��1�u����o�}w1^��o�gx&d�/7 冞��S[օ��*�$�o�}���J+m��1�b���~�`�Q��&k��#W�;O����s����X�tyt�P�2D�DB�Q�ș�p)�R�!ߙv���ZJtc�.����}��4�e����2w�(*1�l�j�['?Px^�h��WD�8�v��qoJ���D��e�IC�g-��'���VثJEVX	8�����d�Mj�e��=/;��R_bK)��u�x��Q\�[W_����u��PόH��m�w�!#dT�}�N�hm�]����¨!��`i��� ��}����{h�9�a3�eHud�u�4�K-@mɩ�����]���I/r��Q��V�tb엑��>*�O>_;tT��̯�.������+mD.�H���i�l�|���a�\{���U઩<���Z��JC��
�py9D��h���=��R�h�_d��_�P*2�e;VE��iڠW]�
C��	�QF���7|h���A_�>�s���m��i�P���s%N�/Ūj�m��h۲b�-�Ώ���t$3B��v�q�z��w�H7	�By�y1�i��v�S������ߺ>֟�Җ��Bm��gx�I��$�|~L�{�[R�e�G��J�������^Jo%�J~V~Fi�����������������j�vU�+R�����v�k��/�	�0x�{<�!
M���T;��t����P�6�+J�6�Il����Y��ρ�h��O1��#/�ݦ<~�H}��^��(9���OɄ�|	��j���P0c��t���4J��ω�#';��s�޾�7&N�ط58�IB~@'O�l��<S�4�N��1����Z ����Jr�� B��DlR��a��`�}i�m¶ַ� �g�!C�d��N�&�����u�t�������[B�|ȷ��6��Lb�t�ַ[�ʀ��c		f	��ϻEfL@N���qx�~"��4�j����k�n$#i�XW�^9���!��M��S)?��RP��(����a�Ύ�*����T�4���7:�e��š�[ܶ�4����FP+���d��{�"�$S��L��3�󿲋�s����g�k������	˦Z�||�ܕ�k�M�7�����?�Tj>�}-��������@����?9k�<\C.O-�X��E��Sc�)�8G>{�x�D�\��u;7�14�N����U	b/���a�)'�q��"�[�?�}����謁Ow�7�lr��i�����G��1�������]����{?ƏL�1���	?��]q�Ͷtω�#��p����(h��:*I�f�W ��3���ښě��݈:��
�$��̿}��k�4�g+G<�������y�_��4�Zz]�y�$� ��Y��Fk�>�Q�-7봃5Ph�Mg(��(�@�G��ݩ& �I��S�Ҭ͠�U]kɒ&�X�W�����Ͳ4�֎7��O�lB�|鼒r�m�]T��M��z���jP�dx���35ǚ��郁{�+�C���L
o��ezC��&�0�z��B�"��}�zi�r9���H����s���EΧ���Nu�B{�rV���4C�,\��.��)9!�[���?.��+��?&�B����w���,MC��f�_˞����<�8 2^�З��S-Y4��[����;Vk�Jl�9�l��Tͦ�z��n5܃�����i�(���B�/�����v���[h����C
���m�1�JGӃ�-�= ��Ԣ��&(	d}��� ��_u��&v�_���F�VDox���^*��_�ER�� 1�8�O��y��+G�>��lpq��ҋ,�۶Y�2<?��>`$������s��[4��eC%e��{�0�m�r*WB^�(Zr�CFk��퐶�=}@��j�ӫk�c/���3b0|�>�7��n����z&@@���5��ڒ���*q��;���e�7%2>!�1M���:�O🸈�|ƶ"ĵ��:�Q���ojV�F�!�Q�m�Xߦ��砎��|E���0����8�Fx�<�6�^�cb"���/�ώ�-8��V_�I)?�rܒ�p��W_/V�.�8���9<�����	ƒ1�����]�:9'u����f�YD�Bo+��wwz�uv��x�_܏����_L�&���L�^ -��Z����D�[�ˈW�	��n3��5��@�n����R�9�����|_�=o�9� �~���+�0z3�=��9m�Y�����K�W�HHb���* x�݊�5��N�(�%��l�{-؏��K�A�rb���v@r�M��c�l�i���_�Ħ���O�Gr�'h܄Q<��h?�I�(� y�X��8@d9���~�/��]C6@�,��ko��A�u?��cUA맆�57�@�y� j.g$"�$� ����q�����Ib�+f ��c���C��̽�?� B^�^�2˯���`ׅsMi �2�����XyFԽL�L�s�g��潓7����)!m�
a���s��|���eNo�*(�m�{;�Ϫ%�?Q�ǭx�g�a{����	=�LHg# ��$4\�^�sc�cѺ�*sgti�*0�A^^�3���Pm���������%���?�n)Uگ������Uku/V���B܅x��@}�ԶWQ���%��ZJ��3�fe�@*�&v��%.�r��]��F�SmH�m��,<�}/���F�-�ukgV���6�Baׯ��U����*��j�]��o(�I��$Z)�����jj)�]���W��z'���]&�ɣ����<Ęj]�8�p�K�SSS"�p������4��V����.I�4�oZ'Se����%�7?�"W���.2����X}xSHƹ�Ъ!Q��;��
�L��F��Z���Z\���N?Ӹ\�J�,�)I+˴�*�4��ſoJ(s��?��V��I������<����B��7��p�A�͟ô�������#$m�
F��g"� �����v����>���������#`�E�xk��+͹�U�%����Y���\���ن����~yY66�MR?p�����V����r�t!TOj��ه�ZoC�وB?�Zo ��?m���q��������l<���DB�S�*��2��B�;!a!bS�-[��(v�Ԕv�VH���5he��k�O�-p�"� i��X���풏���/˟�i�eVؿ.�=�x=3#��ŝsK֊�O�Xu�L4oH���E&l��X����b�*�}����"�Ù٪�GzhS�E	�{+S�ƥ*�1�_̾o$J�=�I�ıE�n���jI�r)�g1'\f��ޜ���@(��
��ɤ�*w�>O�)�-B�'��C��L��ŕ�&3ZY���2�=��$�#ގ��|���y<p}_�3J:S�mEE�x~�Yn�����/]\R�s����ЍMa���&x���4�x�	dR�߰y+�կ#to<�1���L��S�j�������
�ﵖZ�iFr:I��G�����Z:��P �["�����{;q�%��A��"������)w��%�h��̎%��k�:13F&e�m��>�tBnn��qiԖ�ƍ�P��g.������UUL ��i??b�g3� �*��qfw��1�ٽ]�����
dx�E�C�O#��D���		��1J�+�a��Նq�L9���rx����bRի3t�Gژt��
�����N����6~�� g 軳sF���.�:ߗ�xN��[�dM����@�>|��;l��Z*��}�V�R86R�ȇ=r,[�J+s1���~]�d9�{��V-��㞠�+V�S�D���'��3Y���>�e�������k���,�T�p&xf�oȬMı���ætAoL)�e`0G(�����c����j���뎽��� �4�����^ws����=�d(+��Mē���+�n��M _ȿ�u"��g'�ʗS���V�l�p�k[r/�iA"���1��Ϭ��o.���Y���(�	�R��4cc� ��iPP��45�o�[�B*A2B#	�t�� �gs0�PAD���:n�j�:2)Ll��q.��/Lk�fR��;3�3�������*�zO����c���.�ߙ�e�n��{2oMH�n���^'�'��8���[�l�z�3��Z��4�-�$?��P�ޢ��Ym�s�-�n/�z3��pi[��k��@W�����������)e7���u�Lr� ����ǣ\H[)�K#�9��%���m��W��
��Ñ�m��Kb9��˸e�bJ��K�qIBJ&�r��VG%��ilf\>Re�mKX)D���oS�W��1���MF^x~}�V�k�h�x�`���E��I�T�Pl����{l��br��կ[\k'��;�h�&�ۓ��\-���ĺ����#3Y�·��kߪd�q&p�ff<���O�͏���3`wtB��lEG�"[Y�/��p[��4�}+.��	����҆���TȰDE���y�� ����O�8yl(C7�e�/��(�l��/�/�Ko��L[h�aK�]8�=��7�^%�o!bx���챲�H z	6���q��O������y�}^܌�[��L��E^ฎl�νļ=��9� ���L]��=�^���J���+�&�����f��hY�%�n=gRP��	'�vc������1��b=@F˓�;��'
�};����$�*f_��y�֍���&�~jvˡ�o���ml�&:��� �.q�g�s`�Y���K�o�掉��s���..?	":^�석{��%�>F�N)��1����	����|O&�Rqd�D}��9�V��3W6�1�;�������F����G�\����Yƍ��l]������P4f3?)��T��z�����ƪ��m������;�Hxy��W�e����<���d���g�z����Ŀ[�"fDj8Q�g�=�X�	�����`�mfh�����^�v �_1�@�Ǆ@s����&���S"�r��� �>ٶ�*nw��i��|��������-c*� F���ý�*f�1���)j�Z��u#��i�l�����I��	���)z�\��ޭ0��b�(�|��w����w}�,��,�Epl��w]u�tj� >"�޲HB*no�_ ��۟!�o_۱�43md�8��#����Xկ�4����;�v�{mcY�a#�M@ek��O��ʴ���b��)�L	I3�N��Ģ�Ed�3���))�:�؊0d)�L�mV���6�m����2��cآ�V����*�'��Ɍ�ꏈ\�#˸t��6"`�s\��D��x~���+g�<h���HԻoj|���J�0@�[�,s�j�Dtíy���B۸�m�pLV��{�[�3���/h>�&�2M��/!�>�|^#4�YqsJ�[T�TX�� tgh_[q���S�EE���N��_�P�Vn�&z��~��Z>�$?o?m�lO8:t�#}���2㏀E��T�@��F�'F�R3�eXJ�@MߟY�W joJ/lr�J>�/h0���>�g��|��#h�r���9�e�Qlrz�Ι�j v@�AN�P���=U�jc(S�}k���NJrϩ� �cG�/|��Ouԩ��I�'�E���DqLD�$�����Ü՟�C�B���=x֒�K�堟	r����s�Z�cɷ�#�aPxy�@�5+'�?h/N4�c2j�"��H��k:F��N�i���J��>_k�p��A�T�]���wW=� .-<P�L�%Wa�	И+��}6��ǂ��g��*�9��?�5β=J|���7�蜋MH4�]f�Ԫth���$*��*%��W�1��A���3~��(���Oެq�=��R�51�)�y>¼LY�q�K�U�$�K���^�*+Y\�e�*	s��|*5�6=� ��^%��6o]��؍���aOsy�boRB�F@�e����B��$��~�����0��+�H>?��8U�yA3���˓� L;�xn���r琟��s�.�3���"��1^̸rriu�A��w��l�	�A+To�c��c�;҃������]9����%_�V�^�|&��p���#l�w��k$�?ܓ�[���!m���X�rj��#0�X��|���Bˢ�ëMF�!ι�s�ܨ¿��]a�.��B�\��{��44�&�����l���|�]0��Jrؑ����$c�rz��D.�MB��

�6T	�����1Y�3_��� ���K�F�ŝ�}N�R��~�jQ^�&&�-8�|����K���N)�omo�>��-��G��X$ob��@�`����n=�}=y)�=�j"���A%���//*F���pC6_�N��yPf��X���'1�}�3S~�w׿��5�����g��T�\�[���_�+6K�|��"�b��U|�B�����?�~�
�/l;�o�|�-h�D�H>��*L/�)\F� i����x���\͈D���xzs^;3s��r�G�)Y����K�+$�/Q�!�p������}q���9-M��Kk�c��sG�i�}_i��v	]/�G̏��L~�(� �h��W��:�Ϛ��\�(�8��r���#�$���4�04�%av�cZ��jq�?�k���ͧ3�9̫i��g�Ԥ�Ot��-�߰��|L�]�!i˗�v��gēe�[I����;�����n�Ph?���w��f�bE+�y��ch�����9�!7Rv#�yW�.����P$}t$q-hN�QFu�,�p��f�U���jnFѵ�ٺ{���o�4�}[{_����%�-6��1�]0P����N�c,�߽Iv���?�_^L��@�:%����'t�w�?~	<;��_�`Ys�
x��ӓ�h�O(-I]��i{OO��K96�;+��sVX���@�Ǣ4��7gc���:�@�'������f�l�Y��w��.nLv�?�s���6A����� 4����</&h}��3�5z�h���i;����V�mQ �S���u�y����Y�;���jE����ư̿�������{��b/�w��[t�̀�xb�?h�)~t��+���N�N�a�g2�l�ڥN9�҈b�(|�MФ����la{�������eIY���Y����T�%�;7Ь>%�~?�3-ϗ�v���2�=�HH։��2g�P��p����F�r�Ys���3�̉�3�����f=��E��z<�V5q�*X{s�L������W��2����5�q��D��r='02|>� �ڈcP����V�	�]�
���T�z��ޭHQA{�'m�4���&+�c>�n��(;Xp������1�v�m�iIH"4�	�9����}R�����a���;�?�'H/u��(�R�ꬲ��d�p�>���3TM�X>4���g��U\ⶳ-dhO3H�N���(sl��<����~ ��k�:Q�E��G)��`O�b��H�XIP�H�f�:���~���Ox>�9�OQ����Y����K����o�_���r��6�� ��K�mZf���xq��:�o4��gd�i��pD~����;i���{�u0N��=Zy�[V,
�"� 2u�R$8�������N|~�Fr��G�0��ar�A���5�|�<#�2D�ͬ�LL������f.���Y)o�{�ڊ���;c���XQ."���LЪ7��߾8U�_��G����]Y�Dc��D8�׵���VY�Z��K�Y�A��X�R_�;�>j�K��VT|_�m���H9��y�J�!�L�\���7k�ݫE��ۢ�b��;?�J�0����\��ۖ"�\���N��{ypd�nx���h��3�yJ5Eg�)��VN����{X�_���3k��<?L��w(e�BD���S�]<�cZE�Jo�:��jC��Z&���x>�Z�����ǣA?r�Ի� /�6�ԁ�,m�������_�̱հ��� M	��� ��G_�M2����+�J������e����ڎKe�k��Y:��@*KT�\g/�7k���6F�;��*+�777׹o��ԩ888؃@� P������TIR�U�d]++����oz�C=��I���_�WL��Y	� R�f�n��~��wTK�������(�yH@%w}�W�/�����SWL���?����~�.`���ݱ�Z���-&,�6�'��5'�)�o���)�Z���ȑ��t4��r�"2X������"۠ʬ4�����`m{gG����0�t�D��ۆ�b���|�@��/�_���{��O���f���)��Q\�M��=h�y�'�*��K��7O��Bt3č�Д'y���JFC�Qj��H4;R��L&�ԭ��H�k��+��Rg���_6JJ�R#�0#�X&�}�r���}��ƵJH8~�AN���CCC��W��;��m�p�q��,�ƺg��o!xg@~w�H�A�c�r]DkE�wZ��³�zE#3��[����~V�#X��4R����۴�oe(�*���������ǡR��s6�R��߁lg���_rs���߾�'ƕ&J>�gv;�[/��Med���������R�L{Z��bNC����6�#��{�^�L\��z�qn����\C��F�߂9MV�"��[�L�ڊIH�dJ��+�GSEl��ٝq��7��'&
��I)o���bt���՝�$M�6��8���&=Y+�>R(bS��ȧ�U���EC9�	f�O(t/�r�|!?�f0z4C�b!���)��啭���ܱ6���D��� �2���-s%�"�b��-%-u�}��fN(B���a�J�͠�L˻dMkj���'[I���jΒ{fy���f����A���|I�×cL�
�W���bf.=�2���L��ܞ0��8�� |�=�Om���u$$��ú�n� =�۰P%��mN��� �������Llvƾ���6_ؔ�����;�cƻ�Y%��Xd���i�1��A��IB��"�d��</��_���cF��>����+�g�i��uN�;SG)��;M�����O�	�w�5ݷj�����|�	�R1+�5����C:��:����HE8�� w^��$�]Mn������H�������<]j#ݕ�yac���,�,?,���
�����h�j��P ��ŝF����*<��7��$`� ��77q�@_�I�k���� ~�f���aQ|�EGfYEnv�y���w���;c��E
p��(�U��!Ov
=[�q\��#t��&祐,_��?�0Q�[�,P�!TAٰO��\P\�L8�E�в�)�ʘi
�^��^���]���i'�dm�f���*t��2&C�~{�m/bT�HP=>f�����U�<�h7�1�P�R.U�5��>�*'ҝ�J����3큁sk���0m�W;��}�����f��_�ո-^~e�X}�1r�v�K��c�|�2�����ϜӁ6K��W~���[ِ�C���5�{�x�T�@gy��V&{:MF�Y��	5@�Fgy����5��\k���o�R�Y�6{ �:�^6w�+$���t 
��N��*8.�p#%�,Y����zB�o=\{��,�g	A\
����R����_�X�tೲ����V�e~#�f8p�.�^j��c�6I(|����͹�w( ��i�w�g7?���Qv�evY�@,��r4�S{3T����c.�JJ��S�L�f�� 0p�4l	]�����$v����lbf���&?q��vN��$C��2cw
�#k
��6x��:�UT�б7Rq���47����S�~e�����״I��0K{n2.�Q��<?5&�!�J{E��dd/�c��Y'nb��k!��~��v���-u�P���Rއ.B���W}b�E�]�8W�8��^1��#��7/�@	-!!���5^k~�!vq��7�SZ �s���"�?F5-A-_�[�^�gZhz��4�M�9f*��"�P��J��g�X�Q�;���ĥ|������*Ͱ�і�M������]�eJ�q�\G��80���ӟ��H-����RSS�%��xf�Yh}��b��N�m�U���0C9���;��U�m���ڸV�5�p5��5��������0N}�A�*;������8�������)fg�+h.�����2|W�(�|Y����<�g�P%;��R�
[�p�����������;^d/Z<�H�,6WD�ͧ�>�~�K�uZFƸȰL~;�>��j=�Vp�@,�fJ�`��c��{�e��׆t` Y��o�6x|���ܳ瘷���:��	O�\�(��W&���ې�>��q�n�,����/�u>yG��y!i$a���٠�j���!K"?0�O���?3����%Of<f�W��y!o�
T5q�K���p�X�= ����|TW$���A�������أ��|���t����Ψ�s�˰��k��uH����V�d�:�����n��0ú���l�4TS�,U�5%�5nB{i�
Gg�R�tR�`	N٧���m+3b��i�a?���ݢe� ���~��_<���ɔE���aͭ�����&�81�IU����8+�
�c�ȵ�H��h��Rn
��=�,��:{����z��?���}Lhl��m�0��-�r(T��<6*Q6o-��c���@#c[��oO��~q�*��������S��Ui
s�?���Vl)c��Ǥy���w��Y}���ċ�����ew�3��e�7����R/{���D=�۬��㬭*BO��y��9NhpKW�:�f��?5�rq x��p�m��Ż��#���E���i0�~���A��q:7�Ct���,�l�&�����d2y�5���WO�k��c����o�zE?���9�O=�(fƼޕ�#9��x��]�/�GÃ>sIE���t��\�<�ǳ��Ke����(������@
��eU7�Q�0�H&�5�)]�o�g���t�[q���@��E����Y������ѻ���1pU��(:樔GO�#���)j^����Osp��/��k�:ں�� 	r�g�l玌���A-��9���k̡(7YG���k��5��6�1�ZT��&�˛��>$��i	�~���7���2��U9HI�<Γ>y��H_+7V;,�~������z07�Q\�߱b뤖c"�lb�o)�Wg���Ò)J��+���0>�3��&>��+����K~ʗM1��ù����n6v�p�Mf,���r�4́��U�Ù~yeR�_[W�S�ŝ'4[B@څ��"}���������/,"7�].�m��,t���X�:X7G�]��^#�76�'�1M��Z�I���TyU�zn�C!���x��9���'N�H���gq����7BZ�R�[~	����"�� UC0'�O�r7���;�,�x�<���c98�/�r����O���fV�r���S��!N)?��`�'<�cX�@K[���/�2I���vB�8@��K(`#�������s��<�(\���'�EjoVE	ک�O3(�YS2\�����?�ҙ�ҳǣ�ۙ�A\
5���syƌ7(���d�,r�ʰ��E�cH@PiJ�;�Z �����Zv�cwVcw�-�#ئ#V�� T�Y�A�E�ak=�>�Оr`��Y��aZ��!��[�i;t�N��"���)� �c�r�oZ/��1�z��wC���Rp�c�^�.���ڦ?Y�%o��Zj������+Q8ʟ�}�`��P�^eE����0�����[@@ ��㉻/���ys��~tq4M3aX��s�"���U-��J�#��Ƭ�E@��^��,�r2�4������Fa2p�~ᡩ���\���qUYYy���-g0]�ۜ�r�s�Y����]�M�K��Н7�i{�sÛ놬f�㨀�-akc�j�Q�c�z�n���J���ٰ���	z֜YĄ��7wn�� (�/�P�������t-�~����u��;��.X�	�$9�E4;��c��n�[>Q>=]�f
W�ݎ�,�'�Γ���8��t�����1������;�9H�Þ��da]�sY�y)I}�6z�?B�%��������]�Wks�����1MW0��1 c8U�䣉�3�l'ƍ`��L�X�b����z�em�+2�n�-&=� =���ɠ�m�-�r��Lm{�4�D����ҏShK���O��M��f��T~�*�9��U�=����y�&��p�4?��/���e���l,������g��ڳ,�6e���VP��d�of>��g���S��o�O�T�KZw��Yx�����az���3�`,e���"���+��|z9��^��k��,� }�{� ���hP�Jύ֚%ͤF:�E�j�q������,��)��3ulz�����������F�/�^�/�p���5R�r�����Q���r����<Sסp�ʦ�)�Ԗ32�D�v���m�, z���π��J\1d��fj���<��ڨF�;�adDXk<Bw~[&vc{�w�ۄ@M���o�qpx���w���ښ����d�4�AV%�L3��I�)a�ih��OX����&�J���p��'��}�-��o��5��>Mop/�\�&��|�mՓ8M4�9�{��*V����<;�A�U�<[7�����S�ǖ��̡'�a�-b�n��M\uL�l��F9+��!���ǫe�UH���Y�aZ�7�T�Nao���.ޘ2OyO�Kw�3�R�5ͅ��.���IO}!U.9�FZ��17%�=�������,�� c������u~�����W�H�
֝��[V�lC���V߲��ɡP�V��q���e�ǝ`�L��S���g�tu;ٶ�9d�t	4��=��G�xܯ)�yم~u���<H3��?����m�0�Ur����@�����#�öK~��֤$rG��,�:y�_������ ֣&o�ң����~m�x&�K|_�*����f���s�X�X�Ywm��]��i<S���O�&��CE*o�X���x�l�/L( ^�&���1�p��8#�S,�l��qo�u�Ot��M]\��4��jeV=m��9�T�����[��~���R�rxV��{�/����y��t�L��u׻�]ކ�#���n������?�����@co}��N�O���[n�,��+<?�5�<S˅����Q�2gۥ�B��}��{ukV�����7��>��v}�Y��B�aM �y��ܮ�8��'\#q��hq6�a�E����%�Jp��C5�P�=����qq3#����TN�����u������=��	��f�]���n��ƨ��&t���.��㌷㞺kU���)�R�n�>�6��F�߫7lm�+�xϣ���7���Z�����[��C<�O��<�7y����(C��'dni���I��3�W��e<X{�M���yx��q�q��1�^N��U�U�<A: ��K�,�v�uJjj�n9�b���0�����5T��q3%r^S��j�1�i�����]zɧD#Wxx�{i�&���_&k���QL|
���i�Au7�nf\:?����7N=�2F��2Ř㜍��v�����,�����m��}ZT�%�+�K����/������w����'(���!��追��tS,A�Ҟ;�.֝�ܹ���5���"6KpSJ��Y6+{��Բ����5C N*ך��x��ڢ�F��1VIS�B|%�rZ�n��!�{;��P��m*���� /t:��26��8�͵�*��'W���=~�u��̧#�=I~�t<~�^�^�\B^{8�5��Ű���8����{���*��ۀ�����[��Rfւ��BY�z����?�}��P�G��g�7	�P�zr&c:2�����Y��V;e������!'a���ϫ�N��tb�,a�5�u����t�x�ݶ� '�-�������C�i�k6�I��4t|�m�*@�����.�r\>Lp5�0=õ�L�:�(�p\�6��A��î{YU����_�x��͔��-�ž
Y�=mp���~^�î�}s�\�cQ�ٳ�������q�J6�R�,X���{�o��&�£�V��#�Cr%㖕5��� m���T�j+d����?%k���?I���C��d66��x2���f�)֘=��L��ϦB@u�>}�"�Q���vC
�����ʚ�n�pB7V�3Z@�y������<h �@ō��ʉ�
���P�X�a .�8`�w�.�XA�����H��ǖ�4!��1��(����Q&�PB����|�`�K�;��gw��נ��-/�G9ٶ^*ޜ��N����#�<h �q��s/��ϟY��^�O�ޗ�4Uf�Ou	�8k�*�LM��,���+����X��0�h��0��ؑ�:��>Z��]���Y����!��U<��j>\��x�?Pm�S0[�M�1g�On7P�5	�w4
��Mb��I;���*���n3�Ά[����mN�N�J�������V���qZ+��}am�] �mi:@�M�Է��ThY�r�L��c���g%Ir�_����b�+X7~�PvJ�k|�#߽!��a�>m3>�<�ۆ���cn�V��O�$O*��=����6G�`�恉c\3���ɚ�S/�G}�ǯ�F
���]�	�����|v����^���\������&h�H�J�ox�U�v�l\�A^e=">�A�mH�$�<�i�5�}�wL[��B5��
�8�^ �K���w�ʤ��:���S�[�:+Bհ}k��= ��U6�i�ъ����Q3TVM}5�%�z��O�K�!�j~Er�{��mp�5q>`	Kwe�g��g���b�����,��OD3�=�Ҵ,u�D'?XLT���@?�zw`�5ͬ-�W�A��a��_J�������]Ǻ���L�~_�I��)����i��ֿ�1��/~��r
�����{ul�m�V���>�I����,5����*�O��&k������`��w��L8��e�����
���ȿ����>}M�h{�?#'اrɇ��W3�����
]��Z��Ms�E�N�c)����S���ק��*����R`��ǇQ���V��N�M�)!�����OVټ+Mm��2��BP�)���@�ؼ�B+�$(��z}��Y�vV�0��."K3����Yߩ��~([�,)pU��,�(\����1���,��ۏD&ݙ����R�C>]9;N-�rU�5�"j��;�1�kv{���O�.����8�U���^��vL�U���tS֭�d���
C�22��]�)��y��
��K�K^��&�>/8�����b��^-4�5T�1ȸ���,��U�6��Ń��㐹<�*t�b�ʡ]�eb�������<�,i��p�W{,'���,F}^0�␿>��e����;"��^/hii]�uy�+ך�m�)lmv�7���:�@c�ѥ����|��Bf'��/�3�%K3����L]���e���k�%��"�v�e�R��5]�'#�cx�z�e��S�|��쎒��O`���g��pw)-K��O=�
��n��� �(E��&���7E���Yϵ$��F�>1-���n�y�y�2��7	FN�WUpa>>�T,N.��Һrf��8I|V�)ا�\Q�F�k��G���3�������x��d�-��l���SΧ��g�Q��O������&���$�f��6�x�/K\+E������xrV%�y�q�D�O1�q˒�bD�t�81�N�+�h��!߉ى�3?6���)ei����;��*V��Ff��n|+�����鲹��51����U�R���= e>C���lA��b�܀�₆�?�OF^��Y+&300�YuG7��^'x�k�NYg�������i�$��y�&�d�`)���y	���_)E�+��H��_:k3N�m��k�ٱp�|�\Ф��ǔ��h�oM��������X� �����iW��%����~�m3ݕ''<���g�W�����:��͟����N8L�5 ��r�*M���>��4� ��t�[��܇��AE�mOM�$�S�,,@y�}���Bl��@��<N�a��%���V��/�w��>,�a�&��hk������2Zۆ����%DZ����chD���a�:��������q��9�?�\g]k���JU�?�y�9&ȥU�Pښ�*-�D ;�Bd�$d��J�v�����g�x�
ߡq�wt�{͘��%�{F�ʵ���Lo�,VE���%�����������C���J�w^e�8n0!�ϵ��i��O�n�V��n���;����y�e�HJYѽ�̀����5S�c��O$���G���[�Y���d����R�խ=�>�f�O�m�/z��4�A��!ϧ{>��͕�?ܜ�{����~l�'����{y;h�L�ˎf5��u4�%p
�69ٻ������Wo/)�
9�:F�>�Yڸ�q�z�L�c������Ҡ������*�o��}N%�O{?T"c�#c�FaW����H�V���}���h�k�-=��(`��a|�o�k�t�_gT�O��,}P vQ�p�+(=�ٸ_Le���gRtV+��*˳�vD]K~������4�-Pa8!����������/��k3���t^�2��3!UӮ��������M��gj}���;�T����v����S��x9�ي��w�OC�#�68P��o��󦐪4�G��X4�I�?/�SVcy�c�����C	��1ڼڎF�i����"�t�)�J��U=꩙����O�HcB�O6����^�=����
WCf��Yony��*
1�xC��Ť��Kү��b�yE�+�o���gM']�)�PN�J����^�����������GF��Hǎǫ�a�~]C=�D(Ҫ��,�a �����K��T�i��ҕ;�0%�p��A/�0��?�u��Ms���9g�����[�
�|rj,!|x
�`�ǍV��6\W'T����V��?&�|���]�!fb�:����0{{�Z4H'�����=,s+�6���'�A���N:�Y��<~4���b�@aQ����H�:�CU�{툃��o�$���g6ob�}���Eڸ�{��g/���"o���
a�Un�'J=ɗ�)�3���A^]ǿPx��p;ֿ]��G�|�9d�9i�j��7�M����;')����� ��)LB$�de7���v���lt���.a\�5��q������$0`�r4�~{ᤃ��l\�[r�2vU6�&i�|,�����ȯ�F�:=�m�?�����x�>��{��4�&� ��jo�s�����"͋�FNwF��l��u�=+�S1qY�+dC�$�f_SB�4��u�E��~����4��/lGǳ�c.�`:�>�q�����r���_g�gQoy��U�sI�;28}�v
���������,�F�/�\���s������);쾖?Kfk�y��ZQ���j�x"��C�/�u'�G�� RB�{4{#�[���Q�ͭ����%�ʩ�8��s��������^"�xk+H�\�v�X���N���X��b��.ƞ7n]%dk�#���k?d<���}��I3��k'��}����s�+�iWKN?�Ok�.i��I��(	��Rӱw?�Vh¢q�4����Djp���C��C�g|�@T$^;�$n��>���kM������ok��fρW+#�gbt~�Ǔ�y����y�Q0�b��	b��#�����Xo�]$�n ޖ���L��RE\X��D�(	i��u������dЙ����t��oe��=:�����}s
s/��V�Ju.˯��u4�����:������$����hiAOߓ~QS�Jx�Y��ͲM��8�k*��I#\244<��;m�=T���q��zc�v<�m�ے�M�r�������NZ��PSq��Nr�����n�>�F�(I�`c��R�)���gaZ4�Y�D��8t���в=0�$er�p��,G'[x����@�ֿ��RH�놕�M9��Lc���=�ݘd" ?��Q��`m��n�U!��|��x=��*�$�瞇ү.I�ʽ[�I���5���5���s�8��s!�V���Ե�J� ;�5��U�*�!K#1;��[s+�\�[݆�p kMN����䎏��~���~��3���H&<�=����B�*-Q��\~��xk�sr�ق����Y�0�ywY)n�9���R�����C�G�:T�9��l��5,��[Ѯ^�^}<7q�k�@j�
�U�]�.�w��4Ɖc:��-(=l<pi�~����b�'A��	�DL;�����װ�QLL���&'E���o7�e�܅b���74��(~�8c^�'����@[�yN(��,=J�/�K� �� �/5��J�7�0ˇ��;, a�����m� 3}�1�։�ܚ�Q-�ޙ
;��ϑ<�ݏ!������K"u�LXZV!  ��(|��縒Х���hC��jW���*6iJq�[�.L�w�d
�1�n���a�r��Ϻ���/�ey� ��2ǜpX��0�.�!�n�y;�|F,\A��)��>���4F�x%%�"��>�&�L=z:�w���JM1�n����m�~�����M����-ⲁ�K+���1�++<"W�	�Φ�qA�O��Lb���ZY1a7�]��@ ��ɤ�4�pɵvrR���M���WCQ���H�hz|���>� ��%n<����+��:y���7ee�^�ZS��Є�Up�,��3֗ QI�I	�1�>t�>A�������>�s��n�5�v��-����@3wQ�p�g�����+�^f�Ѣ�d)v��QC�S��-D�O��I�0ON��-���_*J^V^}5i�N�ɩ�z��s� ��:@`�:�?)o��+�Q��� ��i3^�e+_`�"��6T徯����D/:�7A�������(�{��#� 4�������_mm4��Ʃ�6�,j��D,���W���(�� �"�n��6r�P9���_*�/����f�)s����m(���aM�\�M����E�(�A��֎����L�`���SD	�航����.�h�Ƥ����e%�Fa;N�oP��0�_�&&��\�&��1��8�[�@3�nF�{#j܀G���s|lj����?�(߭:�q��ыF�ef�Ч�@i-�� ��N\ϯ#��}}����EOHT��;��0��b��ܜ�xF��bH��T3&y���՜+�1Q�ΒrT�ؠؼ�B���s���xc0���xYV�+��bO�Z҇��X���P%S�`�P�?�B����mBڞ�T������xX���y�׿t2:�_WFM�l�'w���o�D���H�/��#��qv����N}�OT}Qu�T)�,!2��]�(�I��0g�>�ݳ�g��Oy��xٹFz�B3a��{�:Γ�g�V#"W����w'��"Oo�$�5���Nf��1�Ӿ�T&'��]c��m�Ej���6��p2g��hFA��d�����l	��0W�k,3Q"t�~��Z�+SX� �~�-�#� ��<����r�F��+�\�����|���3K\܊�
�g�RE�X,�2I�$y;��]�zS���朋�.�v�i�G�9�_Ŝbf��y��Y���u���3�CܯE8�����V�TV��-gj����S�fc��T��9~��~��G"4ΥK?�8��@ �y��R�6�]���g�^~^�G��~��9���qTl�{��C�!5�̏�v�*dR,��<�H=�w����{̗�0$>� (�T�;�S�般:���Ws^w��S<��ү`���HF ߟ�>���V����l�]����\��@�â�}#����\��5�Z���5�~���'¯�&��se���J�b�ܬ��,������U���) Si�杘��Q�ms	�/xq�^�&b�;y;uz�]b����zGt���@i��\�^?W��ERt��㩂�7t����מ�鎋k䕴�V���VF�Հ�L��^�I�U� {�1�Je��ˍj��=_:��\`�yN�o�x��W�fSo*�,�����4��T��&lU�M�W��D��x} ^��,v�����~x�u^���M���fU�$�)0�����h�Q��7���jă�z�����0��* 䗗�@�Й5r���*�Q�éW�Lh���4��&S�i��ǫ�)��o�!�;�'�1z��$���=�)v"��V�J�����z�V7_@gk5�+�Ƨ�Ϭ5��71"���\G�_u$'��b��]t��8&8˒�<�Ͳ�KJ{c ����"�Y�_0�D�)�n]A���+�&�+,6�����v���+i�\���8���'~zGAdǥ_�+
��C  ������a�����8�w���@"!�|�Շ/�>�����


h�x����1��@`�����K��n��Ӧ�#�M�3<K�^s����)4k��������<<����~��MA�oO���&މ�'w��۶崂��_�%�#<j��"טr3-J�C��x�"_���(�r��n��]�T��(B�)�K�_1��[����- ]z�+�;S�<����T��x�?@~����6�%�GF}�����X��|+h�yE����.[!P�YNy�!wCh">���9��@��]E�CK��E�m�'=$t� n�ӡ�pr��������x/x�>}�?����H@�J%��ٖb�����I�uDY�������o�T1��dZQQ��}����ζ֍�&�M�����z@��ژ��
c�l�����L�!H�n��R��#殞8O�]��-�l�̘���٧C��Y�1i`h���-h��s�2��UZ}@������U�v�K��Z9��څ-j��6JN�[���o�	����*�-K_��~��Q6NR*��"��o٨!��ڪ|��K�rO_������F��;Yj���y3�?�ƸH��@�2�'N����6�Q:����^�����x�J�f0��C�r�n��l�l	
�������[�Ҋ�X>#�8���F���s	�mN�w�,�!�Ζ�}!e�1����A��&���:�y���L�m�_T����N��|3��g��h2�߻]�9�~����G�z���t��$��(�x:-��&G��L�7����Yj��
g�򞉪���[��]���SU^�Eҗ���Z�ۃ�h��&C5�2͢vk��R��_�K�TB|ַ3P7�D��!��;O<��q}9(��r3@�::mE@���^��6p���$|jc6)ca�h9���E��+�Q�F#��]��v�/��<�Y����A�������c�\��~O���j��P	��Wy�js�vǲ�^�±����wdŷ,t��Q�ם�;�/e�(7��m�6!1d9��\�+���p�d^uǕճK��wH�F��ϕMj�'�D���hhp�ڥƩE/JK�tl�CEj��#]�i2]������v�N�+��N]�6=ӛr戓�V#���pXFrϰ��}P�sg�~�'牎��<�2�»F_)�Ϸy�~'Lن��4U��D�A8��E{���q��<�_�O���lmm'y��_m��^\^�-68ؤhB�LT���A������㮴��̠���!>�����]�� k���Q�-l���ypc�I��;�ni�:����X��Ĺ]K��I��&C'��#���I�<Ж�פ˴����Yn�C#c�����,W�rΊ	w�I��3T�r>���/Ge��kKo�=T�m
���5��b�ju\G㚻`DP���y^�g<�����%6���w'j��0Oq��V���Ĵ�|��g�W�t�$�t.���_�#��0�Q��I ))ys�ґ�����F=Y��K`0�尼�E���v�}qW�fa���b��hC��3�9�÷��m[�Ѕ��VT@yj�d?�!x�nQJE���$����nװv��q��7ݷ�.a_��+l�g�7�>�B�{����y�K��ܿyy=5����6F��aۑ���\�y+�笗.K>�o;K�˪>��R�}l/#`2k��Eo&�݉<D����Jk[kc�'])�u/���q띇����7�%��N�[N3�ֲV���M\n`f��5(���+������𚲼����gN�O�Ua��A����.8P(/W�P�X����	�zq}m]���tD�fݦaL9�5�Ay��i`m;`eT����\������3 p!5!�������Y�S# y���U|��A��:^ a%�dn����}�{�� �/�A2W�
R��L�A?Y�'������No �����'� ���aB��i�;I�<R'��q��]Ҳ�EM�)ݼ���;�&�|��}��z4l�)���p:.���q���`���|�"���b�$�%L����!{��\SS��UU�yy�i�ܻ�Vv����\P�C`o��a�DEP|b��e�����w?䑼	�5��֞`3a��:N`��x�u�H�.cGw󇣂ȣ�n���L5��G��W� ș�b��9�pj�p�#�K⢩`�:��<��$ݵoCo��-�,�8'�9��T�D���G����Y��8oweV��9�W�]���䁜��P���+{1�Rg�n���[�U�V�����R�JH�����J|rrrݰkU�ݝ��R3����:����Ȟb�$K)p�1+'3��bh������0�eK�Euyl�x�%鰬 �����[�>�u��_b�v@?<�1f��dH�.̢RK����b�h���	ͤm��Vg���f��1�h����'h	�J5,����"Oĺ�8ҡ���1xSڃ���F���j��W�
2����L�\�'��Q��������ϕ��y"�#���g���l%�۽��W�ڴF�48~V�^;�Eհ�Q^K�G�4��(*/�+�,����Bgm�J,Z����+/�.v�%u�sM�n/�먺��X?�
:yȩ�;9p��@�	U����\˅u
s��1��CܭO<)�ү�����l���`��I"��J���&�G��zG��{���0�q�R������	s
�t�E,��u2rř��~��'.�^���3eaf=��0*��V��]��{��Q�%�#B,��V,����Z�v�gG�a�x�m>_������i�޴6F�rpw�����]���/�x�xpL�&ùF���Ař���oK���A�2M��[՗Lh���A���3�4$�\H%��1"�k</�L]��HZ+t�����y�[<���@�zYD\���8���� f+Q7o�:�<h��X�n�6f�#�V2R�sנ%?o�9�gּ���b!�
 V۠Ôk�VࢻFz��nY͏��_"O�p��f����< ċ�@��O��E�|�����U��1c�Oa�?'/mh�.`s_�\��Ee,�w�g����z����w|�fB���i���~��ax����R>��2&MQ��ƕ���+�ֻ�Rrrg7H�F���׎�y��E���lA��e�֜��2����Zq�#Da�(39j��[|;�S��l��P�(��w�Ǚ��R?]hՙԼ4r3�Kd�^�+KD�t�������r{�!��8����,���Hnj�ғ��h����� 3��Lŉ�w��H�3��~�`k��K��v߳��[���,{DZ/�$'ȴ��N7��}^�#++�H��E�~��#�K^�3���$�k�ʐ_�!��]�;<��L��W������;�&Х���Q"~&(Á�V%2���P�(�ϼ=�	s��n�>`�}�+����d~�M�䉌�.^�&N�T�a��l/�4U`-z�Êz�i��ZGy?�[���v��B.e�V�k��Gs����B9MpMF�l���	��{΍F+���Z���j���E��5��i����7��v������v�)���#a0�U�D飞�q5�
�K�T���$�`�U%5���}���j;�����i��T���6T��-�p��/A|������ǩ��-���=�jk�j򹏖[�ү:
b8�˓�
p��"�5q��|�^L���ȒLx����5��Cl��͊Q͑W�@CR�o�4#�4��_���
@r��* j��]���I@�o��C S}s�>zP�nYګ51Y<}(�_g��W[���I����'�����m+(C�㳟Nv�>��c�t�?e�7�(����{E`��&$88X���G��������eg�����O���[�w�,�B?1l�i�G���k�Je���h��w�`>	���Q�G�\�c�~#��9A�C���nf�@�0�\� ��g ɬC��J�#�ט,��8�@�Ӷ���q�i.eΫ�YVZ�������l��zɷDkԊY'&}!a�c�MCk�x�ƈf�"�x����-��n�yDp�ގ6�Pe����Qk��l�� �y�&��� bi�´$߶������?�`�7�\/((h�a3?Yi���Uy���)2�$P�}E:��=�eR/X#���N�4yo`}҂�\�{�@�;��@�tݩ�b�6�^�0���)⁇
{���29�&�ߧ:�F#(�Zp�vF�;5�h:*�Z��Cdmדm����W����r�G�85��ſ�G�%g�]�njڕ/q�l��,���E���� 4��1�8�:�ܖ���@
T3�,�qGR��ppp�^�z5؈��fy�y�.ԜY�1��{y�<��גr�d�S��3�X\j��hs�I��I�%`�ώu�0��}"Z`��aǀ�+}�ž:�����CǭtҮ���z����G`9j=�}��4��%!xZ�����Z�e�@v�+�s��G�i��JX₇f�LbEz����U�<ә^ON����7,�X�g��b7n� cD<Qd+ RW�%`[�M��1�kt�[�h���U��\mYƊ�yK��ˊ�bRy`�U��ܨ��%_�Lj�/E�����5Gr��ǈq1_v ��Y'k��Ϣ��K���ٕ�P�ﯭ���k
�R֧_Ϻ�Go�U�HIt�������N4f~�5Ln1��C�d�.C���:�GC�֧��w��#a�Y3�E��oM��(��Tʦ,���Leg�*]j(=�H� �N��^�o2�� JH�}[�ކ�lO�H8!����Lk{�®ɑߖ���U8U2tg�X���Ga�6���L��}�Y@��?N���ד�K�s!�vܰva˽t�9����ZcccWМ�Z�+��RӾE��, �NL|ÞT�����F ��ys֟<�S������K���o���L�- ���d������FKr����;8����{� ���m:��tz��{<!����=�]��L�e?�&�'��ʦ�OuW�ڍ$���:�E�쬰1O���B�����9z��Ծ�����ᝡ�� T��Axt��z;CØb�����_�\����6#�k��Y�������n�9<I����D��	���W;P���7&t�<����u��ta����-����Js��9Mk��GtIF�7$��~���h�B���Ǆz���-�M�e��~L����G�9E���,�b$��oN�~�@�)�ad� ɸ�.���[����T65��87� ��9[?@�TvL�>��nq38������h_,�����yKG����y��q"�a�Z��JW���G-�$�".B<�x���"��(�q�j�㗭��O��<��RL�;�;�.��lR4�ɥL�D6��5ioj��^V7(ћ����D�zO�3=����ui�-�7"L��}���s<ĳ���V��-,�����d���JJ ��}S����%cN���[��#�E��d��xd:��l��L�hs���oZ�a� Sߕ_���_N��_��n�!�Q#�D_���i�8�)��zޢ�r8�p7����4��o"P4����^��Ru�&뿹9R�ٴ�O�r4���-		�f�����k3,����l�!Z���(�)����w�w�?$��ɉ0������Q��b
)��?P)ּU�KJ�Cۗ4�0N�&����>=o��?�`��l�w��d�?�u��s����S�X��E�c�+R�%R/�R�7Z�R:��˫�'�����K�pk���Y��tU��C
i�
{! ���+ާ�ermpK�����E�����
GY9(HU�����2����+��t<�.��sɞ/ԟ�.g�����������9���"Nz�	�S�M��
�[��jA,�b��Ud-KR�V�q�y�̎)�n��`�U$x~�p^�\�=�?	���_ iFD(���2���{���#1}�k�~����m���s2V���c;U:us�P���B'Ɇ�@0���Ds�G7r�$h�8��%x���p�fW�E�R/�Rꜞ���+���i� �c��j*���h�I��a��ᚿ��I(1�3�%^m5��4%w�wt%��/�(�j��X�(x�ۤZ�?iM�/X;8�e�����J�I�I�**�3�ړ�|����S���z���g�l�N�fnO�InPQU�GZ�l�#YX� �4�!u�C@� �� � p����),FĄ��
2�暺���g������j�"}⋳c\2���s�뼻��Q��9ћ�7�7���0�J�Hơ���4�>��q��#n�9�*��+��B��!�'����[\F��q�m� �o}7(�J,[aC�_�ՙh��S���l˦ꪅ�,�	��$��,&g��j����[�:O���^t�.}���M�M��հ8�%b�7/ۯ����^�u,r� ���X�8|r�	�pߑD�7��p�Y�+F-ᅏ'y�ϭ)@���5��xNB�ۮ�R�˂D��E|���}�F�!?�jG n:ռt2���CkV����KM�N���x�,Q�y ,f `��:�v+$����.��uz�^ۀ��b���*�
����E��!}��/���b�觺@�h�͈�7	X�d0��w	A����}vT�IE�UR�"ؓ�	�#)M7�h��>s�Ya<���]�w0wi�fp�.�fׂ��?�ym���o׌��=e���t��'U���Յ��n���2�D��������M�eO�X.'�m��'�H�nqG�t�0�����վ<��I�f;#i6)k����s?�	H������|����WdA��1)n�h�v��X�N1�|������TTqޞЅp$��������T�B?i.q�""�?*�s���!� ���`lM�M�}�7:w2��h�ˤ�&����s����C�;���I�@��c��A�_ʖ6U)��rE�5�l��!ݎGB���P�����R���?l�AS	���M5E
�V�fң9�A�G� ~f������o�il�	��ʬ`�sf�w+ �w�F�F�w~�B���E��4��~(���<�,�_$���Q�#@.s�9�p��TUU�o��M�V��&��D��i�9��hLf�x��r���N�>��K9���_��߿HĹwGA�]=��F��R��?K�{��Wy!%3�����Sf�C*��vwzu0�S��KG��Xh)5O^j]	7%�q��j���C��A�X�H���x�߮u�o3K�z.�=h'�����B��POe �80�S(PE��d\�E����
2U��3s��w[�E����hN"�f?Ju�jn�XTvv&�gސ���P�Zn��S���g���I���=g��;�������eNo�?�6Nx������6g��/��4�K���pU����A��~G�"�9�#��e�1�Q}�����$>���o&��M�>��O��K���n�gw̷'�1��-Z���@�r	˩�:w�g��nt`�hv�^�Q�\2� M�!zfV�\�J)YK��*���FH����_W��c�5y���Ǻ�O�k��o��0����}�|la��4r��NtLG?m	IT2��ܻ̽7s��kt8]�1��P@YlC����h,I�ƻ���z�3��>z)Xo�n&:u�;"9�����������iGN���D��G�J���
C�͜pe��i�a9��D2`��+8�k���e�ECV�W=�TѓXՁ!�����?ֽi[ZZ&y,�?�gKz��9�U�)�3��?���3����b���֭��{�lzr o��À�ȵ��Er��B�*oء<�0���~����b�Ԓsq6鲛�We0����f�"J.�	.έZ�*�[V㠛�8,�t����n�V�ρ���`\��E��>��ֳ�FJ�}ܨ����}R	���݂ՏZ$1&Wx&�D3�G�ٚ�O�}/�u�o~�3�％�,��.D��: �e9�g���&X��s�&��WyϬ��t��4L�q��޿�ߵ"G���v�<W���.u}/�������������oT#{��M�z5P:�n|'	"9����?���8F�8�����tv"�ZM3��\������a������%	u�R�6)-��2�[^X�a�f������A�:s,��S�[��lG����k���Dq;��,xRSyf�Q�����C�n��p���?��H�):��<9� &�I�J�1��@���Y©F�"��H��}��Π��Q���B��]q�Ӑȕ�XJ%�Ӽ�T���ت��=-��EȔxd8>x��|뗦ο�qބ/Lu�pr_w��utG̻��пO�q7m��%k�فxTr~~���}������P���q&־[R�g�>m��ێ���_��-tZ��WԢ�LP�ԗ����h6_�����^j�k'S����s�"��<k/�/l�M��*��l�.0Uj>�0ѳ^���:���
i�AÄ���(�nY��]�'x{P zȻ�|t�ΰ�#�5b-f>DF�e���ʑb�eaq�y+���u{6��W�U�N�S�{x���eJ������ĨKJF-�:���r�N
�I�U;(����Vm����"H�U�̲J�ߍ��U��z��H�*�½����h�.��#Ű�^�����V�|�N۔�/�R_��yEY�h=���P��;nG���N�����E���Kf�_\\_�&����~"f��-#i���=�}||`�Hx�����,xlL��n*��b�}h?i��ť��J9w~N�y~2-x����m=��������K&r�a�m�3\��E����!�fFlt��T$���!�c����l�$s"����T,.2v��T�+,��Bt�l����Uخ�*�yA�S����6h�!݆c6:��N����T�8~qR���s�X /�ֿ^'#�8F1�b�]�B%���sጉ5p��Ǜ-�������W2x����l�	�Bf�&w���M+����r����f�'Ϳ��Y�<���Z�/������y�=\mއ��:3��C-,�k{��0�dy�&ؽ�W�l��M��dXu�?s�|UY+�~�F�pA~CX^d�d��?�i|�q2ƒ�K�ڰ�0��pMScC?{I)�a�ӵ�T� ��m�x��O��gϨ����y4�+-ⒻL]�t�#�f��7�k��w^��Z|
�Z�e�ծ=j�c�a>Ԏ9�錡� n�����:Nen.�4ĞP�%p~�e�Ap��rq�nY���C}�m���;o�Aź��tǙA�Dv.�����D�\�^R������z!�`2�M�tL��q�,���:����䧏?a�Nnd��V�w��
���/ �;��J�z��I���(�鉏&����{�)bB�5�����2�֑�6p�oS�4�H@�y�
�B��L���yOu�����
pjո�![Z��7�\�T�c��h1�ؔ�e:&LYj��dp� c�i��G�6�qMn�-�V��!��;�@LĠ���t��gC �Q���Џ�dl5�����N�E�Y[6�fX��3|��,�W/�[�y�W�����0{�æ�?f��T���������A���� �E�+�r\�j�U)���Лɔ�w�
��S<]�M�جM��t�{
s5_��b�VW �݉,ǳ���*�@ "���\�� ���	��FF5k�q{�p)th���>���&���p%l2V'�Z�9/��>���p���Gڣo��W2��3�2|����us�j�"m<;��⭄��.ڟ�`0Ե�uF��E>O���YK0�M�u��a�-,���c�^^+^	�C��w}z���q���gk�`�X�|��]�K{&|]�F�$%0�S��t�+�����[��rZ^)�������ۥ���'+m7w���1�>�εV_��S���>��z��;�7v_�g�����V�m&Hg)d_�3��wi�==�1����������;[�"��k?)�j���Ύ�ׄ7ՙ(Ů�y��/�RBa1��]��6f���XJɨ���S��h59D�Jʨq䃌*R�VzH ��-��Ր��iJ�tr�s��:˲��r���(D~�>�e�I���Jq�]��l�_�����6_ z{㜃T��K"��{��5�W=�7�nP$T�sB"���U�l�%^��(�2�hTv����c�%7��[�����lEbh�B���XV�K@����[''ޙ
�9��%�����5)�r#�Q!avɗ[�/Õ��;�p�W�&��O>���8�l|%�wk�.��[�V��}8�ɉ��h�?ο�n̝p!��Y�9��8�­�^�F��#�`��ϪDI�����v��P�#��J����G8�_�-A�K����q�@X�D�����f��,��<��H^��gwj5��\&�uC�y�8�Ȟ�yB���\�ׁ�`Y�+���,S�v�{�:�FZYE��e��Ï�\DH�<:����d|��7'�?�����ʂ`]ht��3�̽M�ӝ�Jd{�1i���X������;���^3���q�Iݼ��-VoJ���ʺYڕ�	XG#��0jB��{J�`@/�f�.����4t��M:�R�ŃqT���i�EI���r�ܾ���6`j�D+@º�b9븶�x�4�0�i
p�5�bv���Q#6r�Uh�Bx���O:lp0�m�-XS~Ȟ���ʹ�/�s0g�&��~H�a���Gq�zh3<��X��N��^�̯]���k����H�O#,{�\b�dہ|�S�@������j����~�����W�_�\��9r���v�=����������94�i72��/]���i;����t��r��w��M��R� �E|`�V(���8�x	Ε�f!d��VQ�f����a6�d�)7%�\j[���TH{Z����7}`��k�k��p���]�Y�w�6��������0����=*���o
lC�T���'��"\Kw��O��}�S{+_Q�L���˲>����� 1Wm0���h�I�9]��K�zv�
3��3
�Tx����\�5w]V�:}�Q����[�߹���="j��v��)�8ߖ�W\���X
p>p��h�0�ZG����x]��-)1.++������:��F[[[ ���=��y���Vy׵����O�v?�@R=�Pu�;*���5S��`��B�B�/V��O��QuM��ݰaʎ�۫��Y5Ĉ^(0�hm�<&6Q쟎_�z��G�yb�.�-H]?��wZZd���ű߹��@�=�zu�T��HCҕ!o��80�����4�Ѫy�*dDk)���_�\��f��GՎ R��R�}�kY����`�s�=�3K�(;�;�IEs�x��Ip�l�޲M�����2�̯q�X��'*��22�Hy��*����� '�[P�3F���4�a�.�������G���Vђ 2�6�L�4I_�1�g������w�x����]/G��1�_M�lD����A�!X.S�4i�$���o�lÓ(���~
ϩ�n�!�T��n&�C;�3&��8�q�7c��J'J��f�C���*���'�(�r(��֙h�����l�T��Y��a�,�m�jm�������=�K���-{L���3�r�^�ʀ��+��M1n��>fc�?�F�m�?�v�zHҦ�:G�H��G5��w%�JFOV���&��e{�$:�NbU����w?i��h�������0Zd����q;6� ��IE��բ�SC~4��X����Ug�@�.]�&r���):��@h��|\���r�FQ� ��ۀA:;��
	
o����m&i�G��5��Y;K8��W c6����'
:{�jd*�+�.�H���6'�h�,�p����z�|���R�@�7tc��P6o�qGA���U�A$��!}�J~�
��Z_��ob�Z�C�߮Rc�<Ē9s)AWs���Gr��ީ7��ZO��'���,��þ���̓[�J�sH��z����=7���^���V�k,|,�7xv �����!���D���T�
�?�VI ��m�V{_��yu*PT'���lI�B��>�	��v�/7c�vK�"���P;W�6֠������cY+++[���K�K.�,�f��"�-�Y���1Y��6��P��,N��<X]U�^�&(V�C��O��e�u��Vz��ă6���&f�Ku���_�m1��.�2�CEt[r����T�A�H\�Dڿ9�����?0�+k�cP����_D��� �H�" �!�!"]ҹ"���"-% ��� ��H	,]K�ұ������=�[�qv�3󝙏�sw-mW�=��|jG�O���V���¿��ZN�ۦ�=�=��[�۬��!K���	�������t<A�o���XX�;"wKn 1�7�	]�k�=2%w?�P	z[�6/�-[�A�e�l������'x(�	W�S1�~���~Ǒ��_���	��-Dh#�I=�,P��ڝ���M ���K��#��b�����sB΅)P��5�����E�1 �%���<n!��2�,�q�c9��W	zV$k+=D�ݨ���E���-6��'״�y_-7��ꏐ��fu}qu:����1=`c�U[��8�Rַ���֩�ǒ��s��.���u�-��X��D�}�7�kq{��4�^/& �R:}�
���U8�?�*�dE>�������!WϞ��� uTT��X��nA!�s��);���\=Ǥ*~�T�����;�I~`I�?>�]/_�!@��~?(vzl��`t��0�� ����d�f��er����w�36�-��A�����'�����G��91��D��!a��DX�S�xZ�vu{V�VZ4�n�|�{�1�K�[�7#�#!�
-R��P�j��ɾW%@A�c�J�W�п���@ѻ<�%�%���G�R�O~��o�+�نw���?\�)&]�x���Er�8��TF�)�2j���kk��0	Ǔ@ Ժ 5BJ�[�ѿ�����toUh������u�?y�lQ�b�!��es��q��]bo.p�xA��;f�Qj�Nɥ���i�z�)��R��1,�"d��؉3/�_���#�����!߸q[z�6Um0�m<�Z�2�?f_D[�߈�+���_�d>U�6��	��� Z��Y{¨n����9.	�����o��t�~�C�q���i�W�ITǻ&��8�uDA��e�?�,|�?�4j/��3v]����t�,K���D�ReX��a�����Oнkm�SnsK)y���J�T,$�Fٶ4�ԝ��g��5�܈�'��oؗ��Թ��H�
)�,}��S� 𥆮iD��2)������?anm&`� )�8���4�����ᘜITG�Ɯ�q�O,��B�����"ވ���e��S�[*�R[��GٰN�OgO�F�X�G�iFP�۪�z�c>�V��o��D���&LV����
-n���L���ֱa�lKa�2
{��%�����NMX}q�?��f 1��O��f�hV �ɧu�%�'餹2ǃ5���MıCؽk	=2hX8�G�j7�1��k�(|iF=Z�7ĥ�w�������Ės^E~���!��h��X�� ��q�ښ^�^��� oSv�r8���r�i�F�jKH!�t}�]gt������13䵃��n�񃛋�xz ����p�@ą����k$t�����v6������/�g�j�W�����+ou���@!�GK𛼺2��Q�>[�i�%�)�,jN7x�:���������!�>��໮�Eѕ7X8�T�%�\w�1o�ϸ�=����e|_'J:�j��+M��6?c��#��8�֭g���;�aC5�m]�� y_����C�%����ɞLt�Wz�tB��s�ns�|g�W�;f�2~�jS��o�3�F�3�-p���>����a����ك�T��.�N�) _��w΅��Dޕi�����m�*}?i8/+cY�ZʡX�qt�%�؉�/~����� ��������)r�ga���A̳�y-b�������&r��u�+�`_y���w�h�hp�[咽<L~�w4BK+s$��4�"Y]�ݱ�Գ�����a��/��Xpvљ�:+ٖ��Ðǌ�°�V�[��"�f�"ӛ [�ٲ�����>߲���?þ�X�?u�F�/��i�^���ȠԮ1����T6_$Lu����)�[���x/,w�&��tU�kr�[B�NR��i)�h����zW34^�s�[{�ġ�T�y���k��?� ��e�����jA������z�����o�b�Lt�6��C������j��S��:�g�V!�@�5/Ft��ܝje6/��!Q\�=��a'���h�#6]����"^7ƛ''1n��5�V�0��y��u�r�N,�Hv��mP�H�Rt4�.���&�`9ۛ_�*Û"�پ��c~��0ؑ)��|�2�DD�U���B@D[����E�y�M��R�-	�=��ÄǓ��6�TV��r
xT�7���2h�x������;!�<r_�e�7�CL�|��'��H虈K4V̏�E��wW�]M��eS���n������r��؋�so�f������5�H$�æ�#YMsK�CS���Ck�`J'�y�_荊��o#��T��z`]�lj!��Թf��1�W��9Y��&��l��,�
��$���((��q����y��
"��u��zH�[ޠW,#t��0!�D���c:\�P-��-UԬg�����ej)�o�Ι~�ER���s����oʢ�������%�6kf�ڣC
���1#r񻭈ms�����)[�[Ǫp���CK�n�[@�k����x�h��T�p��S�Vя+�B}\~�ѕq�<�v�3���Hk��������p���<d�d��[�~$�V(-��Ȟ
�l���{��%8?����Σ��W�pd��K��:��\��:�Hom�߯��1Y}�.S�҉�?�?%-;fg�8Hf^wf���Q&4iٮ�s)ϴ���Vyo��r%��Ā�ILǬ�{٫܊@��������W�&��|��Z�R������טQ���+�0�4�����[7;vg7�3>�1�� h���j�m=��1�5�R��h��}Q�&�a� � ��D$�j�w��� ͨt��L��W@�Xؾ|�����1���W�� '9�����tc;ZHX�kz��X~��',M	裳�H| Ј��M\;����lV���N��,E&քw.1��r�ҫi8�Cr�95q4V�����V��Zn�3g�k�iV�FL��q������˽:��>����4*M��o�����E-3���hR鹖��5&�fD�0CG~d��֣��"_��[�&�E�w֒�Y��SN"��|�!��;)���y��D�b蒡U^�	 n�R�5��Pc�@��:^��c�ZQ웣n��Yէ�+��J��+ɓǎ�Z1SK������1���\>���5o�7��?-<�\�'�pmU���᭦*z��ΙE4[�c伩��E�����ak[��O�m�/'��tXǪ蹭zY+�}Pȋ�q$oe#����^Ѩx)w}Ѡ�ӂb�e��H "��i�ɋi��T��KO�Z�'��q����G�5VY6<��K֌�a��ͳ��iՒ�C�^�ȱ��w�c	��9p���S~�~���l,�He�wf#����b��'���+eR�j�S ��L7`;��ųU1��z�*�O��'J�a_D���K�	I`v�0wDG����H������pSw:�!mʦN�#�o"UÎ�EV��;����KOJHטu�^2����0/��t�>k}U6���(,��/T�l����W�Iq��~X�ϗZ>�N:>1�h��1M��g����&.�jA"I�T����(����W��y�.�e�Y�-�Mx9�iDt��%H7+#* .Ir3q4 �� �̲0|}�#��A�L��y�m�MG�Y���Ij���p���>!�F�V��r�[�(;M��]� �	4@�[c��⦧��)l4Ĳ@CR.X���qRׁ
 �4I��RFu#��fL7��|gwML�v6�h\���f���W��&�6�x2ޭT.N��\(���Az���,>"�����K��~���E�����/�T��������l{�I�	�@��//Ɵ�ހ�c֝������X����1������Xä�L](c���Hu�1�0 ��Q���6�����cx/�C;|�k��yv=�)
���iS�]�~����+�墥��9�J�&x��a�h/$*U�I�>�D7�����P}�x�|8�W��a$���<Q�ٌ��[P�?�G���xC�a&�޾�ɛy��� E��5�=}G[�Ւ�"�u�^�=}!y�?Yq{��)�̅�~t��1��4���Jr5�;?�f��a?t��ܐhd�w5�����!���Y0n+OЖ`k���NCմ�3s4$�A|BL/Z?�xYj�;�Ր�W]hc*q*ݳ� ��C(�����m��0ʵ�-w��/������SE)�\/o�2�$�q�S�ֵ���O�����F��^+l�Y��*�6 '���#1[#?����5����U
W�ߜ)K��)#��^_�Dа�kJwO��
ҭ��-z�7V*�����3�
֠�H��#o���L���n�@��l�����Z��A>_s��>��9��!�a9�c�ޯ����A�I �]CG�%�!.�5���	BoB;�R�c�g-瓪���獪�nD�H�Ǒ�� ��X�6��,���*O:���ps嵙����5�~jN���z��;�O#:��B�=�|�g{��P�.��%���{4o��T��za?r��$H��jCs֊�G�=���Ā�'�V>��E8�P�q+8y�:��@�뵞#�X�^�~��1�m��4)���J��q�� ��M����S�^�,�döe#P�8g�dO~�	�F��G۔5��\I|6�e�� �f��hzL��2t�wja�׹ҳ��n��[PL�$@�d�����W����e��ng��|��7w��Ҿ�y+�����h�=��AN4����C�;;;�:֢i�gg��4p<B�M/1>j�Ư*�9�p�6y�Q$��-�\Qʬ�bl������浌��2oIk�CU��$费��6y�^�H��P���=Nm/�cS���<i~�ν����,��2�'��%lm����j��E�ל���m��+�9��'���v�D�<wN��W�M�U2y���O� ��?[��*%��ӭ�����^`���;��x�/3ц
�3�eEy�o�500�ɓy��!�r5��/p��NV���4�z	U�xߚ���w4p&8ۡ/��d�*�v�C������>�l�ݚQ�^��y�N����Tr|;??_�P���?�s]�P������R��l$������kX���>al��_K�W]��`�/����h.7���S�8��\�F��!�}0��2�i>oC��1���Fs��w��u)��*��&)>o�П�׃]x�����?
��v�x���!,�AUq��m�ZQ~��L��g��\'h�b�e�/	k:�G����[�'�ƈK�����)�7�{�w��&6�3�4��M�?A�'#"y��'$lt���
-�fꚌ�.�ӊ��� �S���9�^4� o��[���؁��0��#�ڒ��{�!n�R�$��1�)�)l���!7-�69IqZ��:�VVR/��������)
J+~9G����9[e�4OI��s����l�Ih�tP���RF桎�ϔ\�g���^`����d�Cȃ��bmnޮ��Gn��qk2��D�Rh!�fZU���-|2�o@�q��t/I�Z]�8��
v��ŭ7P�h�����K�2�W��8S*��7��+*��rS�k�̻�5�'S���f1:�"���d�5z�}�ӫN����$�W{��ƼK�J�s̮�o���b�eBmK9�~HR�t<�׸/�NŎ=20��f�FqAD����X����=�<�T�]���/Y������{�q[����&&$����4����LƄ-��$�kD99X�^N�?^���R�OlR%�u���3�J���7��s3+'\J�6�f�n��.$�Ev�Ŀi]3�l+5���Yd�.�򧴷�(˼�C�Q����� ��z�B���8]�Q��0�Q�������6D�I/XC��X�v�_Xg�m�nJ�5Y���+�K��܆FЖ|aE�w֑R�@��*�m�KFx��t�E�:EQn�x�V�=E&�|�B����M��p���o�_���/�Y\��+&�O%21=����bY}�nk#O2���"���<ޯؾ�0?_�4W>��2��0p_�}��0������ā�U,��o����1�r)�a��s	�8���D�c���F�n_��ژ���
�✪i�%Ne��u���K�0Q���ʤ�\_#�'q�u$�c'�֤��&ӥ~&����v��0�*�����n��H9���g�:�g��pv�[e�O^�Ps���޹��OH��k��v'����߼(A����~Z��z�ş���6�����ʳ!�0wn�b	Km�ڑ�k�G������.|Q��qG���׎u�?��\�	�-aa(UF,yP3_��-ď��>3NhI�f�<��|_Q/������Ў�S^�W�ƆX��!9�=������K�C��h
�c�Tʸ�/+
ό���;Q����Ճ�MQ@���ۍac�s�ؐw̘�"σ(�#�d���\�Z��쒺y�?L��kG�_Zd�&�N6�pt��R����W奋.�扷��<�
:,k��(�����\{���N��ެ�|wݰt
�YȯSh�Å�~t�6�aybA�.2��G��<M�.WC\	[��v��dN�K%�#�p8j���yc5�<�÷��e�����!�3��*����ӕYK��Ye�rX�^�懻$��'d\���._���x�f�P|.+4� ��j7�̍ʮ�������n���q�Bv~TA+.f��?&��B��h����������
c�>)(˕�I-l���8&�a��'ς��6�g�J�*x�<�(�������4�~�3�o��^�D��d������<��G��1i����p,�������I֏S����	G���k7���K�����t�wA�v�����ʇ��G��Їųj�&��i���	���v��@OB��3+�[��'��9VG�Oc%�j���A8�8����~�F|?�<���
?��$�(���<�"��:����3�(ݖ�S\�!�T����݈�P&V��^�Mw7�8>��"����io�n�H��k�]�����Sܚ">kf�pdGKv-�'���n��-��]�w�M�21��M=~�HF`�S���!�Iz�!׫�{F������0��0���'[���aG�7�y���ӳ��k˕�K�OŃe<Y����[x���Q�1�kY�f��N�zn��4��=X�0�S�F�)��g������I��uD����hݥ���Y��b��=WI�B��oJ�ZL�:B�1�(l�C�O�3�������JRDw�F�7o�|@��B�2� '���1Zb"򽲿)�A:���9-��ەK��=h������+˒9��P`��o�����8��]?O�p��H��o�����F;GԆ���2Y����ݣLtNoE�Xa�N^SBF�?��G�U#��3��X����߹�b���w饒s��e�˒x�!�yv9z�7Fm5����Њ��Y��4���Z��ȷ�0�_���*2	tU����(�ڹ
[�^IrB	�v�����La���.���O2�j��5Dկ�d7�n�z���(�L@O�O�_Z"�f�㒸���_�QMIS����)�V�͵���o" �����Z	�Q�V�b���[r%Ha�|n��{��;.�U�9׮�i�A���J�4"��/��G���p���vhBXʃEzr->�P�Ah�y�^�)��Ũ�Wu�P���bE�ҕ=����U���X��80qߺ]�W�e�5����-�5�ţ�hDX2]���$�=�o���E���(�>�,|��W�A;��:+;a�V@���8:ʧ�<�Q��A����F{K❗u^!�H� y���������b���q�1ek&�Q܃���:�MmP�(��HpXGB4؛�ζ�����+�XXLO�'�_���
��{��*�\���I�G��$��\Q�K<5�0t�,�:�/@�ar�C�}��q���37","��T�8����x$����T{;���X��3���E���~�6����n4�b;��r�×�6����ζ��"-�3$K=3��$;�`�:��d�L��U��b� 4����!��rl�O@6#k�/��tz��ǌ��^����b��������Mw>�J����&f�CT1�"�u�s ;�8�tPo�.����!�W�a#1Cd�[^nn����SX���'�\^��~��N�T��?O�������T@m�x �53R���<��K!���fkä����{>�Ψaˮ�h�>���J������΅{¬W���tiS����{撶���d#��E��7��V_��E����ް�X�|b���|����f�lj"��U����]]�U�IF^1h`t�F1���ZM�e!�Ipԟ�k��6B硎�!�@��̧:&�crJ��i8��1��L ���^o�]���r>;�^����%��N�2�b��D��*Sf��m2�_I�؏�����N�ŗ`(*�GI��/X���ׅ�7K�*&�w�]:��he��!<����)��\�d�/iLq�~�I�o�>jc���wx��agyZ,�b�x���{A�p(��xu�d``0_**�[��Y�D��������d����.���_���S�+�@��	x�=q0#�"}+mݘx )��J�BQ�H$�����Bk�D�`�����D����VBgA�mv'x�r��3Br~@����~��f*0jw?q��桢�S�:zx�@h�s<����j��&���� '��c:x6(�ABT�4��)��0�,�Uh�~�V������_��em�KJS��\&A�վ������?�V}2Ƭ�7i����6+]��W��*)�D�JϺwa��׵'�}bh��W�����a�sZ�Qgռ}��mo�Z�|��l�s�3�K"?�@"G��!H�d'�/.c�g-��/�)�[f��#d�EE	`�ܻ�x+r��������<d��Q�;1Nq�_�7P6Lx���\�0�|�+�GO��O�W�`d��Y���@#� LS]�,v�����b�t��9�IZ��|��� �v�J��	����b���ox?@�v��:u[?�men4Pa��wٺ�A�~(h�6ۙ�����N���
�`V��r%2���Lf1]��)y?Gx��}�DPn@�=�5�֣���gh�r�dBO�+��@	��=Dnd���GAJ�gK̆B����3�{rm'y�zz��a��/;�vfv5|,���Yy���m�)R\S���Ǘ(�@�>�GѴ�d./�K���/�$S=�؀����a"b�?D�$��+R��A\�7n�ϱ~��^�q��?W
�Jt�Kd�&T�a't\����X�f���Y��s��odH�+��l��@&�r���x�	�:�E&�#�����f[�:$�4Cw�ܚ�����:�[�J:hM��O%��?H<~ם`���VBk�OX,�Q(Zwd��0����|B,��D_�K�u2��._̶l�<9MMB��{oS���'��7�&�H��܎w�>Y�r����L�__�����/�>C�!��a�?>iY}�F�3�>�w�i�o�-��I1�RC ��,gI���� |��(:x��?��	��=be���y����,AY7:�sغ�x�	�H��ژ��w%w���o���r������v��ں�<*�d�/����s[��|�4^g��`+��Q������S���.���l]yW96	�b�Ǖ����!��}���<�^����|����h~��8����}
pbb��&�ևԑ�9K~���j8�-Ol^g����B��Tq��H��uzn���Q��2A�,qF��`2?�	_�bn]N�c
����N�)�JP��2B&��eE�~N_�¸���g�T� ��d]\[l8-jTe��:d��i���PXGX���|��h��|��G=O��xf������[-�I�/	�4��;z9OW�˽��P/�=��t4	K���'ȲH1ݦ�`H�����h7�����_��VO����_fI,I���]��MK�.����Q"+A$�k+���I�~+�>�#�J+�@R��SyL��jj}�nv4@�c;"�\Ph����'�XeO�e�?<t�w��ߙ�K�MW^
M�ѯ|WZ��|FK#�g��kd��;gҵ�+DYik1[<��&�U<�X�J �2�K�3s""!���X��:�g�ځ��PS`�ؖ�硧F>�>h���5���/��_m�<&�Z��q_��6�`���J�䯡�Oh'��or-�'��y�:P��7#�g�$�'��z ;��'���=Y�*����ܴ�yP{��a�Y����vi^�:$k�x�u&�^\ u��U�d�&O�GvEy20�|Ur��Q�?lЗ���o���G�z�-qS�GL͚+(�$?u�f��܌I4vK/�a6󩈔��{���,N��.]m�l�W��b��$/*5�����؁U��K>4y����΋����[�����f�-9��6>���V6�f��_(��J��,�
�zwh7H̾nhz}���QZ��%��2�[��*\ĿQ�n�@"!c��ⓑ!U��ee �>Z��t���I��7)����V��׽S;��صQ��p�v+ʁ[�3���9�{>��y����M���=[+���V�'Jl?
*��M%̆P����H
K���((�~����<����8��d]�i�4�X�Q��\�A���C'�m
{�(�'W|��j�M������pG�	v<��u>KM	�P��',��oɐD����1�A��	��HT�>Mm9���x�����	陋��1����7���Z�j�8��Ua��?�����h\ 7M8»�����ڱ�X�2@0�=|�u�#:}N��#�n6�Po�:\:.��
\�qX$����L�����݁�q!#ugR��q���9���b��G MȀ�D���n���ੑ���t��z���з�K�y$��T��[��dR^��4��	�{G+�5VT�ku��k�T�ReĆ�!��Բ��ʓ?7���OB{���Ax������wt��a�$������ ��*�ܟ(�ٯW�\�C�!W�����`�ۮ㮻�����2q�1���NQW9k*'�&u�����\CŎ��Z щ��-ߪv9+�����a~��˲�uÞ��+�w�+��S��<�/?�b��g�TJ�H�[xK&�o1����)���x'.��I�\��k�kl� ���h�Ê�Q��V�E��ւ�BdH�h?�M�D-2�nqNƗ�C.��i���� ��:1�g?d�l�M&:������3����^�c�|Pa�mH@9��h_�e���=hO�С=��ى������%����1Ĺy�׌=rT�'p�μcWݵ7Fa�SMZ��םD�|���">�=�0������c	�R�-�T��Kn����S�t)�p�;�f@ Z]=p!�v/�a�)�[`B�{�d�0�w�[��[1R�o��'�'�d<R�+��@�~��iOe:S��a���(���*%1�FJ(ߤ���~����	k%Q5�-C40x��cT�Tx/q�pw�X:��fE���z�?�Օۺ�x�S�a��{�=aT���P�L_B�ˆ�E�an��pP��&1�lW3��&�n���������ߘҟ�%׉�_I���}��FN�z.��j�C@�����������A��:�z�㈃cV%�7��e�F^����^	�ZR�*|к�e�g�WÜ�1��Z�Å��+���& "��y�v�X�(^��:ڝ�*�v�����ʣhʮ�nt!Ao�F@�F��O��S�+Y+��ػi�1��_����V0:̒����'Ԭ��$�'M��`<�_Rd�S�ym��mL�iR�Ud�R%/^~�5�<Wܼx��i,m���C�h^�~��9�&Y��?��!�]� ''�'�XK,&�	�=��$`���^�F�t���=ޭ�wl�L�D�]�t�9��osu|�f'�#�Z�}	�i����l��#��ٙ���Ϣ�B�f����m;q*Y���aM9�*���S5�2�_�W�-3�?���.>����B�E�C�,~�|D�md�ڔmhR!���������")����]jM��L��%@��(
ſ�����d���TӋ
�����UO�8�	2ݘ��;�2^�-eY�J�WJ�U���6G˓�T��S�+`�Gx�J�D��SX�ZدF��
(���}Ʊ'x����9hG����a�v]�؟�I{b�cN:�e�KW΍�r��YlP��V����-���R��x�V���g�m��g�˺. �LC����'�1P��4j��Ax���$��������SӉ�ϕ��;ʾ�%m��:	o�)����B��������u�n�CӝrA�������LH�~ʴ��4}yM�p]��Á�"�tS��1��6@�V���ۯF��W9yh�ʯ�Gz�v_a��3+4�zu#f����q�g�o&�;����:�l�Xz��x�����~{n���C�G���A�|�.��ڭ�/5����R��)��$"]"�fŸ?�y��庮l�);~�g��b�.Q�St=_���&�O�B~��SD*ae�E-��z��G��L"�ymC�Z)��a��Jm�Vy��\b�ѯ?�1�M{�{ϑ�E|�HK�{�"���\�����KH�����]u[�jרC c
�.1C�WX,�K��t�gB�}}��Wo�G�i|�
ݓ�X"�F���hvV��A�(�9 �L�#�\]���G���#OQ��W�}��A�{ �/�8h��p����`���Y��j��h�����c�j�m���p��SA��X�����a�q����l�ʲ��?��Ћv�ҙi>ȬJ�|`Gg�����:`=?�+<=`ѓ{���4KV��3�W:���dL�k��,jR��3i�LQ���Ӹۃ�`_&+�D�w���~�ڿbYW/�4���T��´R�e����- �<�o'��Eo�~\6�j~��K�:����YxBᗜ𩬥�;�l�ҕn�ƚg�-O��d�F���T�ŹXt���\�C�L/��^ltAj����
-gE���J�u�v�����[oL�p��8��Z���;eP�:W�͚����}�0������$I����3>���8��4�y�{P<+?�p|"l;½	D���� E�s|D�u�?��W�lU��x�ט=�K 06d�6�$���E	��O�(]$�V��w����D��板%�j��B����طv��z���痣a����\���p�$�{S�a
�^�f '�j�qX�>-4$6%��K���g��
ؿ����.5����
Y�<p�� f��>j��K)��N�����Zu�鮊L:)�}2\e:����"�Hx�
�Oz�1�K��n�	ZP�g� ����f�v̺�?����L.�}��`�&����©�*����i��$����߰Z*�)e���НZ<��r7���h� v=��g���_�˓�����$
��:nҩ��H�NK��C�9?Q�,��f:��c�,�� ��OBQ�5\GVh}�ܳ��e¤���n�f�F��J��
�@CA#�:j�"g.���m��X�p�#Љ�3� ��F5 ������������%�oG�E�^��&�!!���-���I c����7[���~V��&�Uړ*�JQh�T?�8L���}�kJVK�O�n��gM��%�u��$5f���i�a�9���t���l��wG̣����%�f��5�$�(�����g��f��N�~l�E�.����� ~cfy�52V�y��'1v/���_\�~-����Έ'�#)�)YR�����7��o�j���s�q�(�J� ����$-k>�8��Fak��mR�?p:{A$�A
t/"��a�5U��s�;-ʡ]��S�A��H��zy:w�ې7���&�a~���V}1�|W��Owl%����؟Mvb���b�3�X���A��\���ǔ^��%�<����(?�!�k�r���4��v�뀰b�Qm��ok3}ۺ�s��D4�^?��
\�u�D�^�a��Ѡ��'Q�G>ܤQ$,s���5�����=�=�1��}=o�%3N��oCy�M--쬀B
�G}��0�%�\ω�Yom�ٽ��m#��8�����������%v�ի0���iQ>Rg��J��vQ�X�����+J��UȖ��Z�oUf ɥ�$2�o-�U7�6�4� GZ�q��ʐ�[y�"It���I����
�Z�ͼ�<~�R�=�B���*��y�ɝݷ�w��K��3��,�`5�����0����(�u��J��Zjp�k�!���<W��_���1#Q=����t���˛�'y�l�n�a���7��b�͊f��̈́ٗ���]�/;�����%� ���$�N��V�'y�R<"�������f�'.���8�����ê�FW0Q-�Q�6���G|R�F��u�z�7���!�1�M)���F%}�z�W<bS��W~�G��y{�K
��)��#}�j�s�|�j�""����S*]=y���\%��f�!��B�сiVO�j�>[(� �4?��t�j�����A��� nPR,��HF����~I�O��uF���2��^-��l���^�s�ŧ6��	 �7��o+5�s�x����<7d�D,̶�^ׇ�� �ϔn�JnlN��e�7��a��^V-�M� c��r0�L�p�i��:[�$�Ч5��""x�0�Nc���m喫��*A�Z���'���������~�� �P����)�;䓄��{�R��i=���n�k�7C��`@'����8��X���;z�̻Tn2ei�Si�+�4�y�o"����+ڇ?d�|�b�v~�$��-��Fݯ �����N�;��h���,=	%�G���s��1�{�M��s}��ΧZAV��m��;x���l$a�D	w�h�B���50��o�Bo���ҙZ��� [��~�y��h������S)�<�^��9�C�SE#��OP��(�}���b�q\��a������j�{�]�=SI��ajM�W�}M�@�uƾ������_�5��t���p��(���ϩ=I�����o�fo����\��Xչ�<!ݐ�&8M�v䨐K�d[�!�Q��W.��O��OT�w��wv �St�V<@�Ӓw�n�E�x�S�� �P0#�9�q�GX�Y��B焷c�4T�����6��)ah�j�l{�}�ջy�Qo�T�k�'�h&�A��bI�f�;G~m��4l���et_��� i������2��,��������p�9I:Ŵ�O�f�����4%�I,�9��6�Z0Mu��"Lu�w�.'�Oi�a���W��XT�2t��,�*A.߂ǐ&���	a�B�/�݋���*p����.#�6��ʛ]$_������tm��+�K����ª���t&K�-ʃyr_}�nDB���_�G��s�+<e�	k/�5��֣a�������k[f�j@��
��:Qƌj���{�ݹ��H2�����~JD�b@S�c���~�uwԤ!׿vVv��ڎ�М�@�	}k,�����3+���Jj�1�9��&|@������A����W��.q��3�<)"� ���"vHo�t�LSA]Z�HS�zF�2�'�a=�՟Ĝ�҃�)�چÏHw5C3�ܝ����q�xA�=xm(�D_E�pmw�TЅ�極`ˑ���H�[��ϙ�Dvs��&t�C�w�&��-y-b�o+l���+�Y��҈^rT#�ĺ������w����<=))��M���IS��PA?��Un�����S���z��o��*���mlC��|,��_Ȥ�]p��C����Ȅ��bi=</�1�c���]w,уS������O�ʻ{�s��'kUu�|�;>�;�Lo� ����_I5�U
R��v����7��n��W��K�`^���%2Ϳtf��7��@���<ۃ�%&�%U;օ]sMc^�I�}�+��kc{�\h�9	M*T����x�J�N�E_�c�?�]�3�S#hr�0!܍A�/E��KtT�����D�������P��{X����5��@�b/Qs-�Y�g���`�m|��g+�*�Fa�l,��\r���;埊�8*��5��9S�*!���L1�~�D�x�['��n3uV2�l�K�lf;�D��N��;�W�u��X��[t�~T�y������D�e��E�x��W�a�X��ݒQ2�՜'-A�w�
T��c�{��#vم����'�Ť8�1��*o.OA3��<2�`���C��]�t"�=����4�"�Et�+�=��T<ŦA ��>a��"BF8V��pfq���P��`�c�#������Xa�C�RF�*M�p}�D�P:U��+��p����)���v� ����6�w��d�-ſ����j,ތ��[�7W&��fKx��𮞛�FH\\ԝ	d,Z��P\��k�jSA)�L:�vB�F�݅d�
o+�U�W�������[xE�}a�H* ��#"�%=�4�%�HJ7��ݎ���20t��w@�����޵�>��������]tZQIؐ@4��{W� 6�J�9��}�_L�����%�� ����:*��������A���=8'�F~�����R���O��r���Ɖ��8U���^'T ����~"��4��{s
|�'/9 >�<;oV�bFio��Q�<�G�?绩
ֈ����KtʥI�#aC�)����w��|י�u�>�f�n��<�0�����4�1�CF�c�O~�'�o64���#y'���F�2��M�/6��`[�78Z���˭X��{�_�-5qgz��83F?F{ >:e��&�Hϔٷ�.�&�uD�W8�������<�.[���s�#�scG��K��2�����^c�8cu�	6�Z2�&
��
��`*��� �Qf0� ��a�[>^�)e�N�v���YZ=�:w����H![�dU�NtH�$h��g��+���l�s3��+�'�����:�l��N�����7(��J���O�(Z@W�)!�lb`V��Ʋ����� j&�jD�����\��7�2k�͑�ݗ"9��Aρ�[�ߪ������07���\��T�lN���^~�����'�Z^���Sx�0�ۃ��NL|�':�f��t ]j^���ʸ	��W��d�;T?\�ud�L��_0���R*����ΉG$'F�";H��p���9
N���M���(�ʖ���}�N�Qђ$Y����U@O[z�z��]!��a@��Bĳ|<w�!�y�|=i�[|C��⣭��:	s��X؉��WC��<jY�A�6"�4�uMw��$�d��Oqyi��
�Z�(��0�Źݺ.��]�T�e: R���}_ �2�J�6��r�cD4�o��(�t~$x��	y�F2%i���Y,Z�V���K����f�|��9�	d�L������9A�<��(�� �ψ��S�i��.���VL>l5i���]���
ȋV����Y����U�3ޠ�|!�9��f:u`���i��wh�釐�?���H��AZqq���Fl�	&��8VR3AQ����{3�¼�v���S���~yjYGa�q�Q�m�saۈu�8�ĉ[��z2�nT��:^���q ���*?��^�)�PÕ��ViKm��؟yү�k�~s�v�r�#�\b-P�|�$���� � 
"��I�����a^�
9�nx�p���~�O�M�[F٣���7A��AҽZǉw�\̃������"�Hb��A��faԊ@�\dӾe/F�q?1�pF�㥞�\����5�K���=Y����!�x1�E�Rn���
�pHekzy���C3l���8�5OQh.��X� g�+�C"�W|n۔7��+�y���|�8�9&�$2#��/����=m��Kst< ��v{�;�33�fP:�E�<�OwW�����z����m[��ц��>h���e�}���Qt#�-��T-�
��k�=v��"}��F6w�~_�@�_�0b�?�z/!������7Ǫ�`ǝFV4�\�����;?��Kue_z=F{�2U�C�! jD��OX�oH�۰,�"S���]͐�(Vs���Ȏ�o]$ǿ1��ʮv45CLJ��V�^��^XS�֟}��v��yyBzV�������I�E�
[,?�0��"+���&`X���2��CPU�_`���d�M�!s� �;���c�H��6��˞y��.�&�C{D��69���;c���p{�ո���C�A<�T�-��;/���i$���N����˫���b���`k?�}m����}��83ԣ�[)��S�FV:�w��*+'ɗ��&lyl�#�� %3?p��	��4�9�pѰd�D�»�(]�3�f���_/I7ӈ�J�q<�z<��Aq���oC�9Njӌ��۲�o�Ө]��-m�A�F�r�r�=�Cy�.������c��h?1�'b��׬���O��WF�/ńC�ܗ��#��0R}]l���>ϥ�j�򵟟` П��prpg�� Ņ��>��Ҹ7{��w?儵� ��w���:*�;3�հ���ɒy�M���U��+�*D^<6_�y �u�i}#E[�[mKOA��i�Y����Q�U�geV�k.�h���H-���>�4�u�����&���"G�u~���ƅK������]F�>��h�������D�w1�\�+�#�g������]t�-�����x//G�pi�ң��`�f�/%����r8nI���m�ʥ�/�QvP�:rM���֓��%��]	&�]���4q"z�������<� ͓���y���K���P)�M�\>-�U�C�?3b	8&2��F~���
M�2��ZI:*5����'S�1�]��@�y�xቖ=�n݊�~���$6��]���v�.���!�[�?�׆�j7I�U��m�4Q�\9�c��t�*Os[���Aw�'��խ���={=�Y��n;���t�%^�^����E�J/��ŏ�H�K�`���#pO���c�`G>b�l�KA��+�y�/��~§eNv{iB�h�i��b�L}��3@;'u�vBXGq'j��5O�T�Xhn����,���;�GW���4t�|cU�.��e��������;���������9K`P��~.z���܇S1pp������"��8�.>�mJ�lIQ��J+d�;��X�����MF�~���<lt�h�ap���oP'�
�++�y��5�W<zR9�1�uj�,aenE�@�W��i���UMv<�3+8H�Pn�z�T׵QT[h�<�����ˇ���o�K���Z3�/eI����4�=�r�Z�"0����_&ɼ��b��PJ2����=��-9��[��ͭˈ�u=6S������co��ɌT=p����e��0:�5�4�䊡~�e������8��*�J4�����-�͞˯w���g>�~��婀���{�,M'x��B𠪘��|���T�/�e�<�y���'�Y+�Ś�����KMh�`p|��o�G��~J����z�����Za��f=J��x��v6.\��~���]Җ�4�����'q�B��-H���H������%��/l.�o��y�T��7�_�p�5ݙ�u�y[�r�|��A9���r5�ӥ��Y˟�|v}D|9P�O�.}P��X@O��K�T��s����h�O�l�u��Vy��I��������nvYY���DW�Nw��y(���"�WxH�bԣ&��>�S.�0���JG���꽡�r�yI؍��-����CLڪ�׻��e��;�%�ӹ��f]yu_k��� �S�?�S�}��|l��Q8"R[]�`��$��Ua����=C b�\�)?������ګ!_i؞����n��v�ab�-M���s�:����Gp�_�)?�(�	��#lo=)�c.�ؓ
��C�-���k��!=�/ɲ�Dݰ�Zi�de��������h�7�U�$Fs+LK�p�׮%Y�>�<�i�`�W�O'ߖة�f�r��w	�?��}�n��r��uD�N��3񋛇Q5&��l%c^]�~���qĿ3�G�E�-�14U�̋��Kĥ</8��;�\��H�wGL���d����!���=�����B�kﻨ����ca3��Q��G��n@mI���F�iO|��cY���Uv��~?�޷o�=�Rh���ˊƭa�`vR.��|�ÿr�z�1kV�Fc]�v�/��Z��]LQ�m�Υ�ߴތ5e,�m6D������sG��Hy�|�z7�F� i��e>����v��	0�F�ްj�q��t�l�%򦟮��W�<���K(4�Z?�*7����>ר�<��$]�����?q��[	���O�����Ĭm�R��մsC�ݖs`�\w.����O<��3W��TV=1�x�h���[��r3�7;����=h#;�|��Z�B@Z,���[;��T��ƙa=&B���+󢌔�w���[�&���2?v�g�u��)Pf��;�\��HH�A��I����wn}�ͥ�<�w���_~����ר=�DL��5����} k�-���%��6
�����<��7^�aIp!�ŗN�M�Û��׻�C|�9�;ą6sY�^���DG��n�f>�}���&'DC+��e�s�q�>��6r����a�f��+����m
x��B�U]C�]]iŝ�Q���v��y���>�ۻ���ޢ�ö�Q�>�udP5jͤx�,��',IaT,�	O���WzQ:��䞑:���ø7@��#X�d �@�!}"Y�T������}�)��V��u��1��w▝���Q���_}aH�G ���9�\|�!���X����r��F^�i�c-��w�!�q"p#�n0'����{��0��i��W&9g7ǒ�K��Hn�.#8�7\9"��Ȃ���S�0/�.u�o�(�_��<`�r=Y���je�"���w^��@���]V�0��4kHDR�����ݸ���{�<�ѱc׬�A��X(�@�:���xF�7`|;�D�P��2���̧�7��%��C�3��QM1͉q�|���Rv�k\-|��n DVK� 3����S��q�����#]��UAL��0���c9����?xD<�d��b_�Qo�E���|��7/�[�����ڼ6�P����L&�~��'e��-5ֽ��lc�!�y���OiL�}ص�s|"���:tK�]A��x�n��XZ����0��t�d_0z��^E��W�{MB�
)�^���F��o�
���]Ҽu;3<S��e�&�,�n�
���e9��[k{4&#�l�-v@E���a`�I�r=#H�k����e�H��`|� $ѤK��B1I=4����J�T��
<�u>�T��Z8�6��N�_ ���
�҄���Jꌕ�iQ���a�Q���<��J"��2v�>��G��T�ޏ%j5���q/���H?��f�CE��]�[2�zzL��M��\ZN��LHhOP�E�s��c�dT���{��D:eJq�$#���W�D�$��*;ޯ��Z���(��(2ɪ��Q�<	M�{I�jǈ��s��+E��{C�j����ݥ<2�-+��
�l�2�4��W����0�M*Zӓ�П�UK��6���0<�Z;���ΘV�I�ˣ��c{ȩ�T�|I�|.�/��~�#��k�k�+�r��h����$��2��-l�,bd��I.�^0�#���ɖ�J��L����fU=Β/����B�Yl��Ps�g����fj�=H�`�N�:�ᇝ���Od1h_���ɞ8R h��_���9���b��i�I�8HW����|0R'�-]:�!M��5d�(�iI��m*��Kz#�����o��H�
�U���e�����W���r��8�@�Ŷ��E����	�Q��ە�$���/ɺ+�w,���y��t&�I�=6%`}�_@"����y�-�V����\�|�	8��1�)�v��(��I^�>]<I���+�=O�h��ֲ���DH���ۊv�ws��ö.����Ӣ��l�6��y!��7��^��D0�gZ_wE�_-��RN.S�P�EW��oe��������°���M�L`�z{k&���U3W�(�m/�D>*P<�8�V'֘�����/����yC�6������]�e�yXs�_M�^���k.&Jb�2S/IX5�tt���-*�
ܲ
C�D�l�C&��~�+.%�oJ8N�[�
���g��h���_�Z*-��џ ���.��G&�V��-��[,L
���U	x��C��{�S�+,�7���Y�M!}�m���y�~�N�����:�����y��:e*�� j��5b��{��-"k�Gz��C��4���A�w��«�CBR�W���Nj,׀V�-�}bS���8TmD+D�'��(z�����
�N�.�IE`��W��Ɋ�9 ��ؑ��I��W�f�,O~�m��825è@>¡s��-��ֱ:*Q�2�`Ӵ @�����q}�'���!䇈Ta�7���E�~�?�yn���q�Vh��g�\�;��^��DN�d��c߼j��kA�Z^L�G�L0������]p���1�,���Xh�Ρ�v�����mԓ������Ԏ��{C�1mJz�nF�:DEe@�(�q����IǨ���p�۽�e�~�Z�U��׎=���6�!���d1B:.k N�[��+�^H�Z�Q����a�Yu6�\OҔ�}'���Tܯ��Yϗ� �^�ԨX�>s�}��)s�b:�v�݌pf��\���<t��MvM�������%���$uCX�9��k?���<�&YY	���xu�7k|u]ɤ�֗.e��i�� ����^����42d�[SЭ��;<�o&��郺��˨ފ�cd�e���'G��b�X�c���$�r�ku�s���e��y��u��~��~�ֈ�`@��.���pa"0����w�q���1��ix$�:�[����Z���f�o�����OEt��7�D��H!�(�k|a\87�������~�8+�n�n�E�E��*^^�z@���������d�r�"ć�T�I�X�>���=�l�1��G�k9c��^�Yd,4\��ښX;ʧ^�E'����闒�2=q'v-V:jF��;�Y���|䨼Gs2�M�B��r(|q{SZ�J4����auYZ�TP9�+��?��5�u�����|{�����Bq����+˰%�����퍜3�V����|Cim�^���k�s��镛n�b�<Dza�T3�")��Tq�]��
����[�+5��ӭrC�˩��/�|B�#��
��$�+�	I���ߖU@;z�#VN�=�9OJV����)�2�M���j�_�Q:z��d@g���bX�2k脵�W�]W��ep�ا��0���]��Ӻx�P�g��M|x�wLV̓�{�+j0�����vJ�փͿ��ٍGh��Y.6p���.�i���,�GC㕽��:آ�P	<0M�}�a��X�#.V�"��8BkDK�?6� 6�V]�l���T�&��/��h���=�s�����TXIݬ`��[1쳆�T���a஝���V��G�>
�zt�`�g\G��o��7�ʊ�ah}WpK�j|����yS���'=���ɱ�[,H�NW%YF�eke�K	���-!5���	�繖N�h�1��3���*)I��'ަ��W6�����vi��H���W�f~�O�����dv�����lEuj�b̀�.�UqPur�_
ͼ:�^4G��Eu쿶���<�"=H�Ɔ�Ol���~�Ã����v�D;�ja��7�&[o+Uc���Z��xdA���Q��n9?�i�t�\jF~A�[��^Rѯ+n�f��2�e7�|:�Yo2��%{<_��TalP�O$&�N�� ����"i�W [�φ�\�i��.ݕy3�&�P��.K��Zr�� <X�4���P�6��u���#wߙ�6����D��i��;{����_n�'�������%�J���[�y�\���(��?��>�@��b���E�kKa����V[���s���
��cp|��F����OQ듶g���,����96\��	��p6�;om�]@��K�Qq8� �{�)Z��r�5�S������kw >�P�֞���z��Qd�<^KQ���}�<1A܉����Z'y�I[�?ΓU�>�?R�շk��4�ޫE�$ӭN����ME[ C�#5`6�'��� CW�${��[��i=��x@E3��z;wn�%C�HJY�#�������{ �C�M5q��RԀ6B�`3�0	��"|��Q�_lYȊ��E4�]y'��K�H��k�����,����%n/�p��'��{kx|f��/�x�E)��F�cc��4�qȚ9��5��'����r��O*��]6,<<�6��?#���+a)((�,�ov�d�h\���3�N�I�!5�xA^ ��z���T��ϔ�bX���PHc�ue�u�gơ��=��>�а�m��Lb���7��7]�
{���L�����T(KO�t�s�^��N��?*���zR�,�]�������e�����w�N�N��n��-�Zq
�V%}��4_2z����7�B�-��2B1���m����A��N�y���W�μۇ�G[��㝆1�g�Nhph���g�l �㪮.EE37hntFxU���K���#��N�_!wm��WM�>�ƀ�CD/'}Y
���_���&
��|<���hQP�((Ko�!0��x�P���8�D�,���\|sR����L�a�m?�z6k�v(�H�!��=9�2�BJ��z�%�(�)'eG��nj��YA�F�u;����S�f�>Δ�7OQY98b7��Ob����<���1�y�_��?�u���?�%kV�L&���l��^�mM��Q �2Vh[�P�rn��,�T9-�B;i�W��	���Ѓ��[�	D�uԘ���Z�_��5%���"�� #���..bMH��)N6*i��5b��d�����긝-'\S�8��3�˼�BqȘoQܶ���
��?Ca)�ћɎi�wj���M~׏5+�M�꡷5ܞ6�|w3H�}��!�c7��aqR7��>�ٖ�_��7����C�_�+�4V[k1^����C�j&[�Y���#���ѸC�z�.L��<�����Y��h�a�a�����t�JI�su��u�������z~�H �@�ch�ݲ" �|�vI$ٍ���MzG�y����7W�aNb�+�j'1�^��S�Ĝ�r����9��o��VCs.���F2��+).3����g׵�9썌��^�@j�/���K�p�I2%����:�����|���8��,��AU�?m5�ȗ����@+*�)4��PMnk�E�c��5�ߛ��5bѤ���  j�Zc�۷4�#��ff�&Nnq��x�G�dN
c��@ �6�2���?�nf�N^��2�/�(���{�l�3OSsO�x|-����=gd����̐qss緼h�)@�.���5�	�kv����Wx���m���K�zMfVHF��$ŉ�]�_�n_�D�ʵ�=M�FE��r��;C`��ͥ�B��U�[�ʧ�����@i�O�gMY=��ݴ�/�ÁJ�q�I�}X���-��:�=׾}D2���h �D�A�N����m_~vxFWJ}ʓ~����b���!F0}Y��X$?�b�3UQ��?TP������]Bh���p���񓺤g\�c;��lH�-B6S[(�P�;��x<V ������Ps���p��e��뼗i�`��_mI�C�ZC絰�5x�[`W�M�볞��|�������j�<SOga	���Y�E�k��9�s'�"�=�|�#��V�yv��.Z<���A	3f�~�k���=��¡�xH��H�'I�e���;[2��;�m���$HcoG�խ�+��\�����T_9�ayl�X���? �H}>A󹵂��l%1W��(��Oj�,G=I�ZjÀ���]]��A�u��QݼLo��(��M�.y�^%a�?I�ۘKC�ܢ;gD\=X(Ш��Ο���b��{��'�o�Rҡ��-A������f#�;n^���<�~��Fm;*��&������ц!�{f�8��WL�C��3a�O����׸�T��)�վ�Z�%�N�M���i���D�9(�l��f��9v��������X�Ce3_��or�7�+�ʟC[��s���Ở�c�������f��T�	Qg�8-9ݡ��&:vf�k�&�Ɛ���`�E���V�le�e��k�bRgGѲ��B����Ј�ac�nx�^^�Vg�����`�_8��O�#�r�����;�1#��'�v���o�|�G+�&��F�Y�.,%,��������㤆�(\���)�o��$j^��W�7��I��4#Y�tBν��0�XKt�l���Խr<"]~w��^�3�u��<)Y��n�{��F��>����4�[��i��>
T`��8�>T��E���\T|od��I�����&|���Zφ,���;t&�"�uC�m+�ϭ9r���Oԍ���t��)me}�v_-O%���槩��\��R.6�B�j�F���"���rM��;�^� �
��[����jR�	r�zۈ���s�G�\L"�D#�;\�M�d[�n��.�D=	)��f�,�b�" �=�vFQ�IB�Ƞ
�ÿ$��c�~7O6!�&����褵Iڴ������!��p��O�~pív-Y/3��ea�N]��STn��-!A���h^{��h?�Q�R�d& �`Y�	�jk��������Wr��KU^%���n��b66m���5�4��t9.����g�C8�6���d�Nˤ0�R�g�N��b�
��C�(�\(�ޭ8���HG������B��}Y�6��H�ނ|�2<����)�m߁�ܾH��oF�t:]���E��7�]���
�\�rw�*P�$�4��[r9}X��7=���Ы�-��y����a��9�dt���D
 >�3�{����0�7_�@J��TN�-�6,��4�G֞]�	}g��p����Id~��q��&`O0�"Ae�!�|�#A�\p�hB��\~���H-��|*�Vf'Om�N��e��e�>�i?�9��ݳ6V<]�P�7�@�}��FQ��M�g��/�'Q�/r�}�����1 ��S����8�P�u�Ȕg�N�0e�5�? o���ҡA�o����,��<�!���'T�������8G+���V���=A�S1`�٨��ԩ�ʱd�\F��"#/���!�_ڰ8�Zz��3�s}�>|�y�F�f�r���c��gz��V�
~���OE  ����aRjK��7(H�ᔲ��s�H��q{C!,����I�������Z�x�¿�*h��r;@l譋�7�'G�D�{�2�fַ�ć���j���`fe�٨y�q�Ə(훖�t\U��vTR��P��?��s��1��r��U�HnN�
,�����{�uͰ������k�>�z�@e8�|2j��7M�����a4i_j?1^���HҠ\ҚB����[�#��0e ��55	����/���$^8�<��ҕA�t[�����_�[�MGF��v}6�B^Y��xq;�Q(�(lt�wb��#�
�J1�j�α@!,�)5�|�Px��'��\f�W��AE�P̑j�o����$7�D����V:v���h9iO��fA+D��p��f�r}"����,�0�����~=Q
yS�ST�M�V��/yf��"1>m���ѳ\G��H����F����1��/�N��{:������n�$�v��Rם~Y�i&��g��+�����(9��aq�4�?{����$��v*�����g���N���K/o���� �Zj]�8�(?@l���:��a�D�4]&>��sE��Ms�HZ;U�C'A�ژ&���(��J��t�M�CM���"�J�fI�����;�.����fS8^���H�<l{��<(V3�� �i�����-'>�E��P�kf��O*Z�@Mc�<s���L"E�+�K�h�[E�-���vCC*�hqi'�3��]Ɇ�8�p'~�U
�����ˋN�1���m�5E���7�/�%:V|��;8���J`�	ҕ��:��.w^T\T���:*Q�}���-�,����J)k@��H�IJ�x���D{K@�����"�\��{�`�����3B��?i�u"�^�:�+6q2�\�]��3g��%�K�i,�Q��ˎ	���GCi�����u��I'��v��Vhߤ鍅n��@f����F��m뷗B�Q"{�+�*���%���T>�L�ʘ#��~�u��u���B�G��}jG��Osp���nݶ.�aU@ZI�3ܝ2�c���}��&���U�G0�V!�����ħ��7�J�S�����]�"��r<�M�YI�p�:�E-n%V�ͯ�{���r<��g�M|��ԏ̓?���ǌ�2�������G��U`���Z�Z�l{�#�_~uF�{�����j~������N��;�"�����-u��!Of�Wy��3���V���=o!__�3�o��ف�?�+k�]��a822$<�J���6��c�e�K_����&1��_�3��,����1�	��C����Z��*;-�ËaJ�������@z��`G�H�@6�]�7ep8<v"ƈq�YD���X.�KW��$��9?1I�TCQ�e:v����惜���0�]��m�X�p��n m�dH�+��a6�/���>l{fQGC����$,��Z�K����bR��*��@�w'nF)$O�Ъc2�O���xS4ζ'tk���)_;{�÷�C�A����v�ga9�Qt�+�D��qw�
ы�awn�[�S����b2S=�gů�V�7q��o�6�]�,�O�BL�|%nZJYU����-i������/���g�Qԓ��y�::�ꮺj���>;���;g�V�p��G����`��2Zҫ���E�Ya���ƙ������؂%.=܂� dp=�A� i�^�E'� ߝ�Γ��i�Oߝ7t���A?���5��ѪǗ�OHnL���:���1�In`Qps��D/Ğ1߆����6�?��X慎�ݑ]�������.�����HU=���e-���}\ۀ�抗kX"��ԕ�0ֶ����$z5B�+�|o����-Y&aźԳ�� ���z�z2��uW��QHL��/_Z)]��@Nn��E�=up?ؽ��/����k�5Ř7�N�#7�L�f���`����x�:	�v��\]T���￷ P��ne}x�F������� ���>��;��2�_�9�Խ�S�����q��[�l�j�aҬ�:]�a�C���$���2��g�t�B&�5
�)魑-\���q z�X�fȿ��j���cwď�\W#�p��R���I!����|�8�˟�"�x���ˍ��>������S�T�MC�~��
���
.�E���](:�T������׳*�q΁k��N�&�p\�����%���<&�l�)5/-�V~�l��5��i|��\���zF+�C��d���ޮ��x���^��@��H|��X��#|@�d<�����u_~h�ʹ�_s8u��X�o�yu�[R���������֦u�M��v�`��f7�O![ݫ��m�����bk#��'h�C�����J����n92�l��N��#�4�[����_A�����ϙsʟ�8`��J\NuU�f']�&-}Ɂ��b:�����������zN���+�� f (�x�f��D�ןIX6@�mbܲ�� �X��hs�#���i� �(O��9�\�|,�W���
��db_Þz����.�u�G�Gu�����Xf��$f0`�2�^�dw�߁+zެ�� �����;^lܼi�/L����v����=*���P��-�>'�/�fy�3p�e��~hGQx�ǈ�����a*����Id�+J����GjN.Md6c��|SE#˜�	��>i|��V,����!0�������C�j�,���W�3��5y��4A�CA
��h�j\Bc�xB[+֑�\�s�t�Nz�BZ� ���c�V��]�ʿ%Y���V�!���(��8	j�^I��!���!f)���敘��H���%ob\��E�%��^_ڇ:���V��ˊ��C�X���w�v���(aG���N��-��A�+� �W������ϸ���r�MVZ]��G.�M�st�h8tx����%��&��Y(�0w�~����#74',G�����PT e�q�d�kt>�Z����;LKy$#�g���ؙ��yRL�p��zW)��":S��5�X�ل��Ӂo��~��ڠ�^��� �n�X����� R��Q}�� �&����	�k��ݕ��N�(�Iq�d'�C:���M�M�^o��b�L��S�B~��﮲�W	=5�܈07�������DFH����~1�kf�.bx����%r�L��������i$����l���`��������q�S�f�QȖάcB#�|,�.�auh��GmYf�'sƀ��̘޲��VϿu�+��������~	i�jm�,�]�
Ԗ�
��'�߁����٨S���t�j��|��]
֙$H�"�e�A"�.�g���*BGh"w�_�,��p���Q���o���R���A��"ۆ㶋�l`��gP������N܀��0�ҩƇCkE���X��e��?�^�0��s����8�8�T���O��jm���M��pW�����pf�t��r�.�k�%z�"2�C�?����d8J+(1�TQs�w�}�k�+t:�de� ��T\y9��bC����\f�Y�u8c�}t���y�p��IIL�+��^i�^��Q'��H�D{3�����+ɾ�i*z�;��ޜfMVCKO;�q�����_��S��%$
��
q�5T��q���3#H�0�z C�{'���0'b�AZ%��7��9���yVWP�تKhG��IL�`������v(]���qN�T�q����WuD�Gz�k���t�9q�/~B�����4��)E~���j����$��>_�:v�F[jSNj���%'s��}E8�1��0��p1�J(��Z��m���%�����Y��::�0x˭�n�0
�a��� i6F\e�G�U�0��;<��7?iꜬ�|�����Ȍ.��9.*_;g�#�ߓ�����ff����i�j��qcǊ�-(y����'��Q�3~I�S�5u7j�Se�a/����z��XO<Y�$gh#�X���h_4�^��܌�-2}D�jZ��tS��;�j@��&��2���&�7�V�x�Ҟ���DM�Z[��lh��|ۉ�� &ΔP �_p�v}Px��)?S�7z��Y��z	���P��aÊ���.֧-��X�ߑg0XS�~O��}ف����D���������E��Y��v�1��p�vql5��6�5�	Vp�##!!c��G�3�{��kIF:Ϣ�r�Fbd*�ur�{Q9�h�&�?��-g�{�{�ԁ\���'Ea�q"�	b�Eἱ�=�!2�>�B�X��;�B���ⅰ-��' ߝxg�|�����f��Â7��~��`�x���0E��W��4�?���6�8���Mq��ǯH���h�A����l׊�����V�Ƃa�W��k��P�b�M��5Ԗ�F\�鸁���N�(���vx\�V�?�&A�b��R�1k��e���oR�e&�3�m��,ؔ%���Vs̞�65z4�ۄ�ܮ}��<�j�ѯ�@�|���;��5�gϲd���f�6��3QU��9�ʰU��ģx21D����	T�xa��҇�)LhV~Ve��Q.��g�f��<�߹Q dӘ�K}���QiX��xH[=Yj�����?����到��-k�9ŖܪU�]ܚ�=�ϵr��5�j��|��2T1����Lʅ]��t���"U�U#���~�5E�;"��~�jܴ`^Ə����m�њ�-d�mUx�j����si��ف�5To�,��`���%`��Q�u�,���O���lV��1��|R%�t��T�W�/�V�I$��OJcڋLsv�x��D�#X����xK��	��&9Ari��5�[g�Z�ܪC�����+yYՄ����H8����M��p`7FGֶ�1��樨
��υ�YʾH��O2�Q�fY1��Y4�I�x2v��D2�vY�| �Y��5�k2�F��*(�" ��x;��j����>�ۃ���2k8�Ze�Ӱ��,�
����e3n��Q���[O��2��T���G8�������\�L�"������O����ս�^/I�y=�[˄�.��x,���B��C�41����iK/	����&�)^r�u��췥PN���:$p�y����$fGV�̛i����
Y�>\��ۺ|+�Y"����D�뿩�v�UVsȨ��#�ݬ87�Z\�����H�=4t������8l�����ֶ�0�cY~sB<�3����ı_d-���x�)ٯ�A�d�3���F�h�&�ɬ�*���z�F�����@�gl)�C����ܱT�֚��ϙ�c�G�4��V���O�d�+�~ &���/1Ü.������ʷ��x!0��3�L�E<�$�*�&5�=36���t�*d�+'�ٽw}=�8>v!����+Ƃ���g'Zg��1=��v�O��n!���C�� �-����,���o�ц�Չ�>�ptuO��yL
H����OMˋT��9�kd�� O.l�=dkHG{ jUզxt+i� r���Q��ҭ{m�{��������R��Ǿ\iLջb��^6��s�#��p|$p-O%��`��3�tɏ��C8�u�`���ل�uؐ�@s��Z���2z��9o�I6��!�:��X10@�P�'!���ÂN,�\cE�A�w!�k��A}���u)�i�b8[Q��X~���˲�u�	�y�^����g�d��Vws�U}��(����t��+:K�n��*�kXN>712v���:��l6k��u��Y~NK�B����v���T=-vf�p?�����������r�Zz�J�<���\V\�M#�m����Q��F:��V�_˃�=�>1gF��#%L�X^��s�n�@��~����4cs��R�H����h�C(_I�C��'C��m��ez.�XV�4����J�g�k�je��_�ׄ޾m!*"ҥ���t����HJJHF�D�.)���"ݝݱ�	l0���y~���kw\q����t��]N���oI�5fՑ�Y�ӹ^������_�����83<S2"�0�z��_ϣu�h��Ok��K�V��!Y/��gf �8���D"%O�5��k��%&cv�-�y�'E�)aF��b�8hZ�`/��+f��W:h,��#�8-i�����yF$,�C7F������/��;<�[l}]!��)��[5�$�y.�2�]u��{���^�h^�X��v"�+��ǧ�M�V�8�M?�h�b���'O�W,�,��ݷu������x��,!�_

	�~�i�qE[p�x��_N��=݉�I�S�����b�f��h��%�8 ]�z�L�/"^��*u8ZF����(x��囗wh��(��A��n�ܐ- ��I�Ӫ�n��M�?S/�?��c�y�s��Z:b�:�2��Z��3ّ�[��,6ﰖR�m��S�{5X|+��EF=��y_w*�}e�v���[Gc��XX�E�B��L�C���\ԡl����%��z�l���㤘�{����ZO��£ud:G�����'(لpΈW�N�e
 ��_��h�C�.��a���e��I�g��t��kW��g����o�@o�]�o{�M��R�_�x�=+T��'��&�ѼiFF���
_�b�e'���D专p����$�7�������e��.f3-�_$�l��6A>�hצ�����&z=�&|��Yw���9To߼;b�C��#��QM�H'Y�O_��J�<�����[��0
�G�|�������Ț0D/ô�d�~�/�5G�^3�z
R��1�
H����7N#od�Gy�y>U�@�|��"�i�5��yY�䇆qO��~�eQ8�;��r�	s�sR�y+��뽮r׶V����&�:m���I=l�'�-p�nUu,%��f�b	%�uI�/>)O>����{�j�9���a�����c�'�1�9o��H�t��Y��2�>qE+U9���z�r-����@M�O�q�ˎPB[�����l� ��Y#���iGk}�[=b���U��C~ARU�CZ=���&K�h���[����xE���r��$����1u�e �oك�(�j���'�����D6�c���J�l��1����irC8_�N �U-�4�;�f�	˒��p��m�c ����'boŘ�i�f�0O�B5تJ���Hb�aE�;�	z2�?O�5LC�6�:��ɣ�ɔ5]�>`��H�b��r@����O�m�ܳ��W�fW!z.�mx�����u
�C���Otx�����=��v�����l�Y^Ș�Bi��DR�/w�Fi)�$Do�����>tV�y'����590ç(��録����肜�Y/�卂���Y�];�V����O�G��V;�Hd����C)�4;�l	I%Z��Q�qUc�HLa���?�_�e�=Ah���)堋��HK���Ep]�K�5H�Pd<5�;�k�I�J	;;qT�V>�j!��;��}��!��o�c�.����w'C�Am;�h����c�$.����|��1�kxr�C�l~��w]�ֱDkV:��)��x��Z�����慪��m}�z4]������9�5�j�{���dmHOȄ�|$*����ތ�]9͸���"����d2�+ck�I/
xK��A�w�$t}l����f����������n���Cq�7n:	��g�O��=R;�؝�ʹ:Y��1v�|W�T����yx�Z^����xqs�d��-������]j�7#�������S�!��^z%N��j�ٔm���ڥ�H	����?"��G��j#jp跥��2�L�QM�r��Yy>Z����va��Eb�s��9�4��G2d���u��鏭�ą�n����\^�;;�F�}6�t+���E5Z?jTJ�x�`�K)�H:'�(O�.��7y14���Ι�*u�ԣ�W�JX+��L���k7�޿�JA�D�����@�d6��h�`�Wj��b8:Yݶ&/��4�$����gdWy��>��%pV�����\��BF�d	�d�j�r*ҁ��=9BM�s"y�+�L�Ҵ���p':�T�O��8Ɵٸ�)H{�=��=��E���Y��͓��Q��w쬼������4�"[�p �O�VoB���#V<9���rPf�����y�سT�|1?)׬���?��������[uCc|tc�t��K�ŢX����lX�Ω��P":�"���yHL����֍Dje?���0������$�Ug6ٰR�aR�|,�֯t,��ӧE�ku�-���������QN�7��3�����&b�o���x�����h�d� w �2Ր l"�/�H֏�׬܁�F����B���i4S��n���i���������\[�R�y:�H�)������B8�Btwf���>6�K&�譠�jF;l.�������֕�n{��fz+�3��*�����#�۩�\>
 P'��h�Ͻ�s�d<P��(����>6��y��<?��n���翰n/�˓
��ͣY�0��+�)I;ͽ��t�M�����*�J ����ũ!U&K{����
�E�/��K7��*e��e[GGqy�x�Yff�N����͇<z��XU�`�4 ���.�To��v�כ6��]��ZxJ�FK�Ve2��!�>KM���.��2@N2��J[�=�ސ54��r���!����1�
���dɝp���j�=�UH]ޙv''�<�e� �R�O֧��D���-m���v�|��Yg��qVTm�����롌-9�}�n�@����I�ò�7kVH��:����صr_�e|����~!�ו�-+wǄn�]-��3v��E���'_�Ew8����gA�'� ��~�h%�QdK�j7��e�dN�XV4�ޤ��O>8~qE��6I;1�m���5sz��k �.S��r��h���'6dZ�x52LO�Ȫ�K�[�X���3�'�����[}��B�;���x�>���ى,uhfQ?��u~ߏ�&q#���*��j#�;���<�l���7N+9����J�|뫄�bvt^j�Wd�H?
�h��
FF�c��n�<%۰��w#��F;׼s�q�Z���E�UL)Ѳ��ک��L��e+6����C�$�-M(���y��<%�7�����M�qK{V�DVY܈+jH��l�x�䅈���\��L�4�ܻ/x��^_o°o�?�;0�o��c<)�k�3ɑ	�^E�qme��$�k`�Ih:(�J#�V�l�M��7���L�ҩʻl�|fXd�;�Y�&��%�H�p2�a�M����=�|��6Uuϋ�P�����ҋ�s�+S��oE��@<v��\"Sb{q��OܿO�n�ݏ�r?��<�l,;��5'
�2�����6�*���䋌�2���CI���}.)f�9���x���M�`f�4���������2��P�5��������Z�x���"�^�08p�/r/d�E��Ґs1����bff�!I���=�ў��\+�S�g�T�*��˕6ʀG���^klE��.EܧL�(�R~NE�0#�ɕ�Q��A��k�w��V	�<�(j��[-���I7�ɲ��Nu��r����a˨�/b�q��l�/���)�!D<�[��=�Abk��ǜ}���I&iI�v�?�)�;'���s�Q�]6Mh��Tv��'�q�)�}*�T%~���EC,`t�f������&[�B�/�<a�;�;("6���n���!�?�oX<��
��أ��:���ph��c�3o<��_l��^	<�|�������^�5`ڣ�
cj�?��B��=���sG�0vz�q�����.fa�)�y�F��Ot� *��mU�ג�L3ʈW���n(�1y�S�;����7v2�f8�����B�Lbi��ؗ='��Zv+��U��Bz��}��H���o�P�Ҳ����=4͸?o�['�F�L@�J��2�mvh�j�fљ�����:����4q����]}��;&��� n� �k'w��iA7'��U	��`�θ՟���κØ�3�7��J+7�7�>sܸJk7�@-�v	��5k�2S�R6�{Z��{�_t��-�4lk�r��3�|��#r��(�V���E׻k�3�NO���z��I.�?U���嶦Z���zx��ޔ����~��bi}l!_t�Rg���t�c���uZD�Jt_j�dȮ��8�X��Q�m�k~��{e�3��w���:�2�]��Ӡ�쐌QL���Q��$J�v�P���\Nث�욒mP�S�ڏ�s"jN��Hb�LS�x�l;ZF.�I�y��4?3��A������g�9���~�}�w�E������?E����3��@�n9)�V������W��5P��0k�=M��Ԗ�J���}(��brЊ�t�g�A��<�)��;�A`���ؐ��"#¢��p!2�C%{�Ù��ڀ?zL�����2eP5s�y}g=��z�)�c�O�����?aR�"��	�/4�_��z��3�`k�0�;�@-Q��V���|5� ��xN�gG�H��ϙ��3��	�Kh�D�lZ�8G�Cp��`��t�\d<��trh��h���rr�[9C�$c�r�tJ`�6���hU�`�lU$����<���3�Μ_�z���p��Kt8H'�v�<8��6�[�I����֩�H��'K�PK#(�-��]��;bM�E��eg��hVF�G��S��g�MüQ2bIƐKR3j�]�¤O1^4�~���X�"4d:�W��9�r�/�d]�"���/���7�^�t�K�IOt�i!$�L��|.��C4����9�6��5�����]�?{�,r�D�!)��%��΀uǺ��D֬T?Ǚ�#ssc�'f�����M9iܢ1����]%�B�R�)~~�g��W +<��z6͖�JNԨ�ݙ��8�#���ӗ����`(�[��zqlEYk�	Gg��w��ky�wnn�V��?�����hf�pM��,�:��_ժ�4z,�$a�$��euqFH���~�RƯfĒ�������!/�$�LRy�)�p����-��7�k�Cm+?���ޚ����=�2��S�a�ޟcD(���m��z&�!k0�J�=;~l_V������ �|����U^�C�lȆ����@d��\f�Gi�iȋ�"���W��[ӎ9���M)����P݀c޳����>�{+�(V�iɨܰ��iF	��#�����@�d��}�ߒ�3���#s�Oɏ�� Ad8 ?sk����1���2#�-q۩�!����M�C��+��ă~�����%B���5Oh�j���Ƽω����<�z]m�U���e��,�L��8|�+h�9��/cB�/��M�%�Bw�W�=mY!'L,�c:��V�1�Y��i}�EF�5����wm[��ӻljT��!m��ӷf�e�Ǧ^cTLj�x�%�4A�>2�N�ܣN5����7�L$~���D��F��	J���7'�Rlށ�*pӺ}���}�(���`1�n�ɷ���/�	�یr&D~�S��
��[t�� ���6[b$�j�l��珞R��x��%3�k.�,�do�&���L|��g�>�6����z;6���4�~2q�#��>8����c�/�3 ��8�o(��Ȩ��!eu��J�o�w��]���ރ�}�߽�>�m*V�������MD,��%�3:7LX�� B��`�������Eѭ�c�y�ؕ[ѿ��V����C�����<�[��bxNdhOE8�8�׮V��Lg �AG宺�%��§�/C�,�e���M?c�hR�'>w���G��lwC%��;��<|�z4}P�<����*�]t��C�i��>����4O�V��ʤ��E�-��E�|����>ol�:C5��O�e�8j��J��HzlCS���ƿ��cA�/ �a:1#__+} �}&�X�S�D���	@�4�O�̽OL"�3]նb|DP� ��+�
�[�=]d��c>�?,��}<J1]~n���и�'d`�s����ō*J� �ou8]��1������b��m�U�_�8�x�u^OS�*uw��t���'}w�N���kڹ��|tx!����x7"EiF�bX�&��Y�������x߄,Cu#�:R7pHh��hv�� �r0�G����fx)�Y�}D�y�ǎ6rLҵo���Q3�ó���_���9sʨ-����7lV�"��?6S�}�i��	�Jӣ�m�$�:���������j���!�2%z��U��Òxu�˵x���Z}��߃���E�W!9��_�J>p�d<����<��֩^�Hj�j�@��@�@Y5%`��HG@��o$c�ِA���'��k[���;���$��!�h��'�s���a����$�p"<�D�@���X��-!ib8RX���������0��bE�BZVYH�D�mG���$�R7vѢ5;������x� �};f����}�W�Z�]��0G<]$̢C�������ރ������{�H��yP�-3����!D��w�1%S$>a���t�T��`)�� �U��˺Q�5�̯&a8�:��2�6���q���'���
]�i��o���V*��Ђ���E�.�[�@ٍ��-�o
�2�����]?p�(q����ߗ����5d��S����Si#o|�	Y}���y$��Z$q׃)�{�rkQ����۲�>s�%�?Q%�ė�
��@O�'E�kW�[v�@C
b`��]�Ƕ���w�:';k����IT��I� m�Ug'�hچ����5��3ߪ�|D�U�[A�������[���\�ڂn�綨�����k�0�A�}d�"C�}y����B�fvS��
�4~�lm�&$X�>aS�x�j��GKèoN�h�6M�\})B~ ���ƒ6Y�J�j�_`��1"F�7�	��Hn`	6F8�_Ԝ8��B}�ӧ�^�a���,��&�%�>��)L:�¤f7d'W��Ɍ��}!��o��	c����6K���M|d���S>B-���P0G�����2v�ҭ=�4jSi1�d���W,q�&�dV����q��S�Nvp�I6n��@Cr@�������<Y���"��c4�#FlG�^�A7}�)Y��1z~��ڹR�X�t�Ǣ�λc����ԝ=��W�Y�8�*e�e>~푌 z�R1	��׻)G�P2�ƨ�������N�#��!_�O�x�r�	D��]��Պ��N�%�[k0tAUo���� ��6`�{,���5����`�_�W��}CZ�prݴr��ݭ��q:]�
�� �u�"��S�;o�-X�����_��'B[:��\$9G��
���u�F�x%���Z�}8�-�]00�T�J7v��.FB;�A"=�������zc�����OŦ(��o!�z6.�0"���=py
�J�d���Кjj)�)l2Do����/��FC�HNa���vf*>�Sxe8 �U?��ס���/�#���%�'\П��e��u>Y���W~��I���,����'$��~���qu��O���RWw8c�sZj�^�Ԍw!#e���	�ת���u��՟��?s"�W�jciЭ���YP���[�-fO�й��|�61u���-vт<�B5'z}���t\�@�o�@��U�%��//�[so��+�����$��i���X㚠�C�U�x�U���#��c5цg��7e�ň��&�`U5�<�3��>�p�]("Q����c��Q�E����G�7���Y����Ao�@2�<al]�(���䒖�^1_��'eW��`{i7������|�i(if�MAl��<��˂SZ����(���}�K����bG\pJcG��E������6md�K�����&��uC�yR�B��UJ�#E���M|Z?y��� n��vM!i��3�"�!�}�#��[{��{���
��ە�� O��+����r���+JH	��GT�(Z��ؗ>�U�H���-J�3B29F��ȢyP(���l��L�.5(D�<��/�lT�_�D��įzs�_%!�VƝ����s����{�W�3�TmS�Vz��co���kɦG�խH:���	?'b��|}#��r�y�&�4��^7;p�,��m)8#t��l���kkl��r�ؘ? (�ǋ]��b~prrH������уw�k�Mk��ڻ\p���h��2������O��waG5�HJ�伪)�I<�p�p8���O@	��2��w�l���-�g� n��]��̄g!��&�7>L��fpM}D�4�6�.t�,��K0��-�+�ʼb^/?#>�ʛ)ؿʭ�<��gYx�g"ޫH���F�Z}e�� 6d�ƈӚ8VB��f���ҟ��F���-�h�VM_k9̿DH
��HM��O�i�:����3{$*��޶E�E�'`��9�����Q5h����5T6�AZ~��Z��Y�X8NJ��ѳ����ٮ��ʹ����B��g�o[�Q�#�GY�Q�a��(��u��O�L\�>r�����ٕ�8��"S���������L�_{�c��<�����A�=eb�^}�F'���D~>iM�N�CÉ;�-?$���Ђ,l��+�O|T�bdM ��ԕ������Z^F�(��鷥�$1t%�Ǯ�15�ěo��yoe�	!�j�f�	H�i�%�ڬ�+��yB����wOV���#�o?p씱�+�|ҒH-��G����a���5�w��[>������G�z"S��|߇�`ZYg4d��W�����i2�.��&O��oI�ZU�N����X�h6.Y����$��[�Wn����lKl�aΠi���.���S{�\�Ja_����$��	�ܕ��@��s�
[��o<���l@E���!�դvH��nɸ�>��[?����Kk8{�����lid�9�|a���{���t��c׾Ԧ;��,S�7�48�L� :,�#ټ��71�7��zG����}I~���?�]��ԋ �"t�W��� ������&��ETM�^~�D���c�o��B��3gp������SAh+8��'���wg���7�����B���Sm.�@���Ӣ�c���a��8#m/�-��\�aޫ���\Poy�jۗ2�D�L6��P���N��WW��y�WD���:&OQ�'�C͒%�r����s����۔�i���˯�tp��Ҿ&��>����R�}���p1��h�6���l8f�F�z�q�B�|[ܕ�mG-!����]w�K��G҇����}6���d���ګ=�]_���jN�;��@(�i�2�ۘ&�g<EH���w��2�ËKٕ��S~��Jw�ٕ�!�fE�����G�[H�oe�M'����d\N��q�S�ĵ6u�r-��=mo�V\�yџ�T�N����	;p��#}Hzī�V1��)^�&�� �uwl��0�5��1��VEF�w�l�7������&C�3;3�"$�]��^�&ď�ѮzF>�x#2_$9� �q�\5xWy�@,T|����y/���)����)�Uo�S���,����n?�B�Lu�n�����p�^{�ݰ�PEa�b�"Ta�<��8ʣN�v� ��PԮ�%~QEK;'�ٛ�N(�5�E�������H%>t��c���
�-"*�\%;lONҮ�T�d�΁ O���HM%�IMZ�>�&D��w;Xn�M7�Lт1�v�*��Z���G�K_�N��w1ۋ7�C���2�$Ք�g�0�ͯ����O?��b�kK��-�EO�VJ���̖[ٟ:�F��������#(n���,�� 9|��E]�O�Y4»�89ޙ��Ĵ$b�P� up�E�^��r/ ��|ڶ�%Hp�?�(a-3�֋�3x(Y�Ox��vX�Jg�gN-�R�I$uYצ���t����M-��(k5�����oǖ��6̃��#�?� 6�Ix=�`pI�zUZ~�����~\�6D�l�3��)c�J�Νi\"�t�L^a�M��2Z袰?3���ѩ�<ґ�ƽ$y�0��/9S�M��z�+��J�)o|`�Q��m��I������٘����T��<_��;�u!��g�ɠW�t�[N.��x)�qnn�\�=ZD�_`��}��f��V���s��Wt����yf��(1�-�wu�⫽d���##d�ᠠb4ͲI,-�UmJ̩�>a�lsy!��I��ֻ4��S̭�FD����V��%���4�,�ر��(�j�j����0��R�Z�A����]p���s�#�!՜�:�:�d�[��{͖�g�V&7�P2q��a�L��}���ax�Ǵ#hA@h+D :QL[�"Q���D�Hh��!ar����BOO ��R�B�Mu\I9��N2<���?t~�9��˫��v(��J�gp)0��ٔ{,��~H��o寋.o��^�o@"�����p6��v|�.+I�n�w�jn ت�_��󻰷�u_T
oX#�U�-�R�Q�-VX�)�V�g��xYGxN}�o�����$�?���y� (�f<�0�0�~g7l�Q�2�D{���8<@�P�:]/�a&g}�I+/7��Jy�us7ǣΧL�j��~޼��A��dzҩ�OK�F�HYٽ|�9��Fr!1���m#�W���C�i�5ByY��L3}���}���+c��ǲ��l��
{���/�X�WS���&<��2�Ԏ�|C(���SP#��s1�J���_p��O�׶�l]��g������%G<xE��΂�m�'5k�/,�����NSx��B�͞)�=���5� #sƪɓD���\�
{��l�ոBӂ}(�M�St/�7$V���	����hK�͡�Ac��hM��3���:C�%�@���%O���O.Z@]�/��=�}LZ�Q�n�ٯˑ���V�t���[���9�g�̀5���.)���Q���6�ޫ��`�P����!�9i/+N�~�HX�ٍ��>�¨9��[z �R�]���4O)� I�a�,��o &B���H���ϓ��{��g*�����W䑁b���8/���� bӛ3~
�i�,	`|�s$�2�<��`r.�'u�8��Xw��|	#��lOG�fV��/�Ѡ�� L~I��%ԾOy�!�
S���*i65u�c�l���}��J�LmO.��������)����$g5Kd��$7������""��������i�#�7��?���e|�ʌ�V��@�,��uEU�$�qHo�;��������z�`f7�����@���-�M�a@%�ތ}	��j�CC��7Ov�h��l�l�r���n����LS��(Ω��I9Mѥ02��r}J�[�϶��"�ʍ�d.�D�Ɉ��;�b�������^���]WU=C�EL/��g�w�]yi�:,w�������ژ�`<�����>BN��TL���ʏ�9�%!#q�:�z�py+���4��|�u�/�]�$"\�����.��4S�߾k� Θ�^��p+�r������X�t�5*Ư�r�gDx{P���:l7��%���[���2��6{�Z�3.g.�%VQ{�>��[���s\ж�0A�E��{�vj��i����s��\����/�?���d�o���ߎ3	S�-%���j;%,݇�Ps�O�6Q�l/���>��[�D�ڮ��������;��z���˵�����:Nč�h_�Ќ���#t��$�^��4�s�y��w��]��@9���8�ȜW�[�0U�˝GH��f�|b�}��=V��� �t
�G2]�F�%�#ĈV�yd��E�Q��T�a�E:��J�|���f����N.y��8�J���Q6<?�U�C�>�,"��^KX�m��f4��_��*�N�s��˹J*z�6�D1>d�AzƆ�$��oB}CcNtv)�?(�W��3(�_i�NZ�'��Y�� m��ۉ>��e_b�dh�MLܜ(��n'9y�'qǈ� )@�΄��J�.��`a�q���f	��Z �$}�nxC�yБ<O�.i�N�O��fT*y>:��[�x�.��3x������i�������M�Y�=S;)�	��Sǥ��H]�߸�PR+�êll��������[,��jwrSI���^����B��,���rE������K~`_�=�>g4t0��i��M�~'.T6 ))P��]�Ĵ>���\"��ЉX��.ic'\s�32���>i�� �If?����T���_����0���^����� *�~��[N>�<�Ih���p��I��i�f�6ŋ��;J�$*�O���k�@>%���O��<�q��p��-i����+�CQ����ᙈ�!�����<��-G�F��]���=��{׸�2~�-�vs��;���A'|amLmD�
(����"P�}���dx=h���Ȩ�ԯ�xq%���ή�о�N&]�rC����JM;���-��B�	J>2�!">�˛)�M]��iD;2�krt��޵�.No���a_欄nk������6�Ȃߚ-�^��W �a3���*xR��0���ڬ�����@���&�d�&Ո�p|�׊zc�1�VB�0�S���Y8��k�[��=��'���W ��\�!�'�՗I�,ZW�87���;��8�/%�f�>���N7�)"���|[�����FvJ��̩�s��t�\M"a� F��-�+t�~�:����ǨY|�Ⱦ����p����^��Bh���b�ӕwT��d��}Wo�n���aJ4Yds��u��pv�o�;6�c|�o=�|W_�{k��^��X�C_��8�5��ߝs�w~3Dߣ�I�K%U����k�������d�H单Oc�l&b����_Gn���W~�ƪJǧ��p��φ�v��'P��R㊧�E���q}Z�O��oj)��Ie/tO���X:3
�]��D�MZ�b��i���>E�v�4y5YX���<��}{Y�� ~��
�ӯ�N����[��#xݨ�O��f	͓�7]�	Z�0��>�� �Jr�^�\��٘�c1Q'j��=	�����=&����Ϣl�.��'n���q�s�bf(�,��ud�����/>e�%ŗq���s����{�wϠ��Q�z<�6��1�>KW�q׌D(�X?�ht'sGHz_jK��5v �JQN��P彰�,�OҰ�TQ���$����z�tr���jR�B��TY���&]�A�Tj�g� � +&.�.E���<��?�8��3SΑ�l#	\V�g���-��-���!nO�f��	�W��n%����vĽ�}�G@;�V�}v�d�]�Iֺ��6�G��Y�눕��;ܾ�	��6�XV�����ԭtY��ݷ�ӷ�o[�U_�pFK,�w�7���,.��c��-�rK��;����f�Y�K��B���	̓8��{Gg�@�. v״�?�����������t�W��R� �������C��#�XZ4@ԥH"���>��䤹��:QP8�����}\���5f盒7�BF����;��і��V΂s�#�í��tf�ι�ocu������,�zkH������l�$z�q�~C�/�a��̝�i!�Q����Y+[��7��<V�P����!��؇�m���X-��I�)���I�"ƺ$9�F4,���xhX@��q�l�~�;��K��N�� �bP�
ѳ�up�%Ҳ��Z�͗�X���!�P=� �O��Ƞ��>�U۸���ѡ��l>ϑIX�e��bج$��#�<���c��$��n�M)� 8��5��0Ψ�*E*�N�DQ��.>��tzO�G?!?���	�V�;xk`}:��S`u�p���β�*�R���O��i��
�ycTs|Q04�V�yT���	���3h-A �(��.<�+�f��Y���b57N��h�G��kNX�hxJ�\E"jHZaP���k/#)��*$��#�>����D������qq�t$�S�8�}4h?�\�< 2ڂ�se�(�����U{u����LsLn�@�<YJ|`�B=�Yq2z��y�h�`R�C"�/���|���q�
�[3�1�˧�����E� 	�l3���{,*p�DP��u��h�Aws��49+,�D�_o�~M��=�PX֫�	��4;݉�ޥZN5zڞ93�̯*�fВTI�|��I{!R���$�m�R(�~�I]~�(;�-$���'UK7�$��V�0�xe'���ծ��h��H��_*~9$����6Staz�h3���8|�?�Z\"�~t:�#�%�L�~pGZ jؼ�Ι"9��w����R��P8�W#i4��c8&���@�a����u3C�/��D��2Lm̜�΃�,�Jk�#܋�z�&�ȼ6��H҅U���vV�SQD���O��ψM�]U2`�H���p�?ɾ�v�s:C��'1v�.(�q�42��
X��t~U/}�3�9�sB���VƉ�߾a��xE�|��L�g|�)V�����>��R�E�����7F�ZA�8� �V�w�{��MG~��J��F�5������2VG7#�Ѓ�q��I�Kۗ7�+�Df1��Y)Қ��Ph�$��	Ԫ�kB����2��� ep|'l����n��l�B��Oo��h�6qM��[���yI�pv�v{�gk��Gl�K@�Qy3��O�4��9pG�|�c5����Pu���iP��_��ٓ�,��թ��U:�R�������$G3{�b�k.��x{~�P:7\:n���?Ž�(�d�m
��綟�Mi.+�E��?�gb�G���/��*KI话òZ���#���,��%ބM�Smڊ�3�^�9
���v��R飹����=2��Ŗvs'�(��I��gF������g~d��%�a*p�Ӑ�^�;�bh��%��L��$�4骄�+�|����[�*9�v�>�y��dJg�)��堑�t/�(14��a7M\� zԲ%j��8��4p�0���ͼu^=>�i�4��c���[~�)m�q���KF/־��U[�g���c��b�B�@p��$� �وw��:�V�1 �b/��oM��h>���vp����NS��И�#"Pm�S��^�	
�",�g��2x�p�A%<��s�/e�O��yW�Hw�/��w�?OoA���u���|��=��[ �o��.~	�����x%[O�c���*B�ښ$�MW�ı�5��X7��1����Hl��ݤm{����
;�kf1��s2��&�#�������-N�+s�����37�����O�5m
q��ڨ=SL�*I�I�jp�k(�K�1vA~�$�3�]��������Lb{��eF�����)�y�����G�� n�w��j)Et���= �r�ƛ���/na~p�L5���.����8���~�5��75�?�y�4�x4�������u���T��n��y�7v�̴^�B�Ғ�BDJ-��~m�cL/�˕U.�y����mب.Y*�r�/.<�����G�fM;��p;��
���ƥMX���Hbo��4K�͍�j�q(��)�Ia���E�*��6
�%��\����IC%���6;i��W������w���r2�|��->�n(pα]��+|$�KB�*.��HcߵJ[��ޡ��jw���*���'gk�K?�8��#h��ߪ?��9c��P�$��bL��fw@H�b�{�gi&���<�k��YD���Ž$Q�g�d2���$P1��,IIgW���ܴ.�5��;aq��ݶ����	9��@O*L��ΏD���L�t	LJ���n�ȯ!��%xCQ���Ѭ�.]�β�#+^h����d}M]�� ?R�ĆQ�t0�~��b�a3u�r�U�e	Z������e�]zX��n����b=i9�^�ްe��L�E�I���tяʬ�!&ю<�
&Eqo���?�| c�(�îA�o��7�^>���b)�i ��<�X�I8_~�[�.�J���|��ʠɜ6<��|>�Y���7V�+��َ|T�iV�=z�S�F�����j�T�崛��b+7��~z�F}ىwº$O ,�By��3sj�#V�no/��2��j@�o��fM�S�
�gy^����[�TD�/v�!=���
$أ[�\�H��~uhm>0�N���sj7W��0aH1�	a� 7=4-�;������r^>�����ghx6��Y��k��`A���<R��J=�A}��r�ѳ���!�%�ˏ9�9^�:
���	Na,�Z���J߃^��h_vU���#
}��u�.� b��m�>���4/ v\�d���@ +�%��4B���CK�e>?�����zV֤arQ�����}8����X��،�*��_��)���m���,b� �ȟ�9b^��'cu��E>(�?�ӓ���P1��4�,��yG�շB���y,Hj`��)'�֪��l���Z�e����<��	�ޤ[��a-ӊ&ߵ�w.�$�b�j�Us��Z����@�o��R�����ҵJ>vx��/H9������_̇�5��4i]���u	 =r3���O!Гv�zs���H��~a�r�H�ָ����_hU�bF�Q��f9��,i��,Vi1s��g/B�|��_�6�q�wk�'9�xy�g�\��q�bMq2NuO�ɩ�q��Q���`eT,l@�R���u3-��6<ٓ �\��T\�#����m�RU�RiըZU�v[�vmJ�-Fm"�^EQ�.�{o�7�C{�H�������~�{��=�9�s����}�[y/�����M�%���'���t��'�k-��	��Ա=a7��k�kT}�ۛ~��8�Ƭ�����2v���z�k��eMf��To�f�[m3>,k�c��x��&}��-�0q1ٍVk����Iqo"�CÆ��κET���F��;?���:5(a���������~[6h/��!�Tx���#"Jbt� 3TG|�����0|/�0�SRw<i�<�5�L�uTC��_� �L�̔A����y^%\㝙��ݻ[������Q��������յ�;dSs#�k�J%��q�:\���)·J
���W�AE��|��g�w�4M?�Nm�L�찥��T�9��\���Br��w��/@9���uQq�xV q�Ǽ3ܗK�� ���$�et5�vM#����]�
��oT �4�@6ng���l4c��*z(���W���/+�k��gؓ�]~!��1���'z��8��I�\)xEo��6�w@Q����ގ�}/���)!���8��dP
��H}��~�l�����N#�jT����P���hU��0����V��B���{���aB6t�;���#�D���u�]e@���]�(f[pq�^���4=����&@X\mj����u���S%�*{��{o�Bָ`Gna�ȴw%�ؑ�P��G�6'�mZ5~U!����h�6BdǢKzP��տ�XK 8�{�~�5�����OP�r�������wYq��	�N��k�����zJ�9H7
 qaWZ{|vXs�#tď�F�h��B���֓��A=�����P���]������Y�V����K�M3	��)��Ry�)���J.:���2~Xb!�wk
kE��~�c��_.%QƊ��I1@m�TG-��j�nR`����o3KA�K=}?�z�E�|�Pua��!|%o6Q�U��tUi�G��a�:��I�Gɣ��yU�'?�e�*(��+�f���]��܆'����͓�z�y7��
�,�%z��Isr�Kq�s��(Բ��f�N�����ҷ������I�5g�Q�{]��Y����e��ғp�V�P������ѧjlxe��&����:����"ę��ffODF*|Y�X��`��d"�z|�}�=Ƈ���c lv��՝��G���z9�/|�����4r�w���f�
�L���f6�lLA�X�ڤ1��3R�aٻ�d�ڍ��.�{������C��n�&5ayY/o��� !B�{22��g3D�"���s�Xc�}�$>�@��� ��s{t�������A���&��c"aD�Ҵ�(�HʌM�C����]V���4��w�����Fu����}�؆k��l;>��T�,�S�e�bպ}"08���K��38�{S SB�/_��֬�����E�W�h�#�� �������Y����˴�֊�:�o�w|�5O+��*��~��JU�=<��#��*����)=޹: 8��ý}�4.�q�s왮�?��!��jy�G�"*U��-3�9�Cz��3d��
Z65v��"d򳰫T�͟��	�<���=l#N>�Kz��,�>'1�'���I��aU���g�%"�o�#Q:�#�"5��#�=嘼�9z��qNd��Di������_D�]UCw TS(X]N=E�>.Z}����+��֗��p���a �Z�5��q�t�b��CM1����q&�=�^9�dD�쟂m�|1C�Ǯ�J�a��e-ǫ-�̞������'|9��s�ΰ2�F2������P���mS1;�N��ȕ<���!VU��c�������[~��I����_q��Q[�8�@:#h�:G����������|��C����^C2��iV��<qW�MP��I�붸»M�L�9�ބ��f���]���>�(��e�S�6�d���z��-��c��B�"-�n�3z)�֗Sg���;�d�[�/>'~8{4&@�[��>�[�ҽ�q�pt��I'�N�'�pV��-͚�VT&4F_8*ݱ�à�'KODh��s�70~����j���/Iј6�����g%�&���0�fi��7A<���jZ����<���W��ȭ2�L8S������A�%b�g�'qTH�]V�i&h϶S���/|T(m�����>���ϵ�C4*N٤����u[�y_G�[���l��߻P}�ԅ)Bꌱ�U)z2 ���*V/�f6�����_�&h"�+<�!�Tԏ�j9�3zf���el֜���E�[��ǪՋ��2��t��ج��+W)4��$����<��z�ؚk��rX� �bOO�+'��鏻�O9B�P_rB���Q�-��[L��K�K�����k��4`M���2��嘢aMo�q h��c�l�D������lO�طQ��	z^�xR�ݚ|C��(X!a[��������(
M�(.��.a�Ǆ��Z��5��_!siq��@�x?&��;ɉ�p���L�R�{-�q���|oA��KǤ��Z4\��=Jq���~�G-:�f���G���@얱���q� {��K,^�s��?m��ө��r���X��4�J`�-+^�PT��;������M��O�}�}���!�Ƒb�;���K)���p5�y���3�7���p5��f�K�dKM��k�Z��H�^�rL�շi�v��Z.�bq�w��&GGz[���&O4m�WURyB?�UYi�R�(��m��������x+l�Y��5$ ����ûX.7�������Gtew���&�-#�=�<��#�H�cL���S?����(J�)��j�z翆s��Z��5��)ɧ�n͟��&�Sr�cy�*UW���*�L��p�����e�5��"8�{��I�ޝ9��<�N{��e���S'�}���|�W���^�0�*)ʨZ�̉%ؾ�U�c�{$�xU�BX�z�1��޾t��=+��E=��"���?t�L�8|���=�~�3��i�����L|<sO)��_4��,z�cQ7%?�W�#ł@m�v*(�� J�u�_B��n�E��a;�w�H�:�&	[T�T���z6<J}�8������BSG��<Oi��E�:b��T�z��{�r�@ˡE%\W1{d�9�@���(A>6_�ӆS�������Pg(yi�Oʡ�2S�v�DT^`�%j�ۢ�h�Qg�U�W=_�>��۞�z��6|c4�HZbY|�t88K���.�nEⱗ꺲b�Tͧ������(,�3��Ju��푲�vկ���i����w���	g�d'�����`#2�����m�u�K� �������p9�q<4���Ra��) ����O|�2�ձp����J���ns�*���<�7f=y��e�܈�h���g\4�H�e�--�6`�����ᨴ���ٞ?�Z�V�V\L���QTM_D�M�0����@����H��kigIh�A���!vP����ME��fYb��'`�˟"��ֵЖ���:��rً�ߴ6�V�>40�����]RZ�p�a��;�jZD��t���ӲO۶����vjޤ?���L�-$�H��Iĸd�NJ������Owf��C���f
^�'v��_�+���b�^��p<b����1�{Ty��������'�΢$Q�����E=Z;��]�g�v���/?@�#��w��J�.`U���� ��o~��j՝�kx��*í�fw	�>��x���y��ꤥ��)'V��hy�sHe{/�rb����/�R�4_�K��ՅZ�]0}eH��ep�9JBזϫ�=t�P�r����b�B��v����1�7ǏQ>��J�,S�C0�K?�4b���s��K('�"Q�X抌p�jO�8�#�/a�ގ���&d��Q;���R{K��(�$;q&���$�57�Z�'N}ܳ"0�ּ����E�i���܀�ͼKҶT��|�P?9d�'��ER�EDm��N�;c��O}�No�m')���ި�{��魥�l�YiA������36����wN1��0��P��iv�A�\lf�Ǟ�[�J���ؔ/G�.����'���Ӊ�S�2S��uG���?�6�u�Fmy�	����a�� Gd��q)�ձE
c�"�_/���m\߇��������o?'�܄y� ���s�pi�z��,�u���&�	G�<��k�=�ۤf��])c>���u��/q�/��f�
��<����@��/��q� o1r	gD|�d��X����dm��~Q��&Yu��DZ�t{���ֻ2�8P��V�XW$���\�w��cG@���n�^ր��tC��ܕ���E�^#'�w�Ty�n�g;�h�9�0�2S��8Ʈ�Dv҉r}�\�D��-�6s�_Dv<￷��C*~#�� ��4��x�<ظ�[w�J���Y�� �V�9����I�b�X3�K;s�K]Pp})~K?^w"�����~cA�S���t�0+�,X�sd��-8Gm�v�/� ��-	\���%�g�̤+�6Ʒ+ w7���D(v�1t?���1a�[��Q"F����"��-2c&�̻V�߿�>3�a}-ЛBm���ۭ���"��!g�]�E��f��d�eYMo��H��E����E����9�YU����P1�Xׯ�s2����K�
���{h�J)k���t��>�P��X��G�<'83;<��u��y/��<�$|��	��K����MV.���q���j��k~�>��C�]#T��~֎%hkR����$��s�p_&K��PW 5��"a���i���F��b?^����?0�,e����Dq�J��he���ʾH�
.��])EE�mA�S|e��e�T&V�[G��)�~���@Sו.S�ٲ��>b�Al4�7��+���e��L�n��NO�ڭ�G��Sa�$sL=xfi�C��o������0~��i��9:0�ծ�t?�9:�z�z�����=��HF�0�9{��y���x������w��iH�3o�C��w��K(���[��|ۄL��M��w a����ЂR�j�F��^��k����Iť�L���e�&�Vf�uI܁-��_ƞ��N���qKĊ�#^�_fM>����y�c�©ڧ�?	�Q�HFn��x� jF���wA,~����l�Y+ݴ��%4�B���TY�w�RH��_�I�ʚ]q�4bP�A�P�QL�z�w�! ��V����3י�����߉����uWhN�c��\PZ��^�;g���\Qd��Β��
���-H�eYJD���vwQ��t����Q�.6���O��q�[�mC��r}�r���kd,�f��\Ѽ�Wひ��f�|��6��8~^����R_7�!���ґ-=���p>��uA�����Q�7�T���;Ӭh��#aQ�r k:�E�r���\!����F�-�ܞ5���:��I���m+̈N�*��'���>/?�L!)��r�Iˡ5�a��8�=4<gP�tʮMܝ��+q#��7�T�d �(M�z:�4�����H�*c4f����t��
�Nݟ�#I8ˡ"s9ۀPyE`�Le�d{=���ʁ5ړ:�w��\���>.�0fq�Z8�BFm����#����92j�d�����IL�B ݁�����߻�� L��U��#��l�Ǿ �1��]��̧��)���'.��{�O�]?p��;�}<u7I�+w��8m��.U����}�{TG���ϻ��J�*�9�,�t�qy�ZxN,%���9�҄¤���>G�����%=g3\��pyT�@��B�lyZ���'U����D��w)7Z����������VRė�{@��k�����f��O8�
 exM���RSR�i�۸�1!���^�)���?I�w��o�JM��*��/�]�/����(��RѦ����Jz<��`u��X ��&O�h`6GT���.�d��ޱ�3��Ui�K����V��Ӈy b���ŤV*�FH�Y�q�sP�j�co�ؼ��l���?��\z�&KiP��M�j�b�)vyO9�Ͼ�̑��ɖ3?���
_����ңBO����ߺRm*� �>HQk�-���tEg)_�M��8��!k�=��2�@�l$J�z�vھ�P�=t\AD<	c=zb�?��~Dtbd�)�3�L�O�9y>}���-g*��ï8ӂj@d�H�A�ص }_��x�FoU�����ͅӫhp�Ur�g���N�2���%tTS�LitAj�<v<"e]ms��M�������TFH�#Y��;R�����>xP@�Y��c�;��0N�zdm�ڶR���s-��כ��y�8��%�,�ڕ���r�u/��T�wJ%U�_�B��+0�p�!9|���繀䟴��bvg ͑<�5'�"��?Ns���y!���:�]%�ty�$\�����>��; �Ψ�3�u��s�O&�#&����-�`��os�R���ߒfukS�#n��5E�X��-�^i�/�T͢�����=�E�Y��t]���Ol�Or@��=���k~1E(�/��ׯ�F#7^f'��B�^��� �_${bt�8�i���5�����U��xtJ�1[����A�DNG���f,s+����z���|�MtN��d�E%�E�ʙ���
lcX[�Sir��\�@��΄v]���J��Z�.Uf�]���(�\�X�vL��QrY������{�<�@w��tʔķ���O2��"�Z��&�7Ѭ�l1��F��S�ib�8�	���,��ȧ�)m�d:�)��ֿю���mr�ԪJ�5D�����hA���;�p���(�*J�?O
[�>��)pAˑ5-!dУ�ԛ�E2�|'�f��PD^cqNC���YX`�g�����<K^� Ak�iOߧ�v��*9Ĥ1Nl��lmb΋3%�C��1kzV�F�ӎ�^��ؙ��@�3�����}�6�4ԋD��c�Dce�Y�Q�@�G��R�{�/�t	�5�5[d���߼�^)�q �TX�kŀ�w;�[���7ʯs�,⃶�e�N�v#�pe��	��P�� 3�@{MQ���N��ƌNuo����fP�9�"/꣑���~f�Nr뽉\K�Z�{%���f�b
=2>�V�|b)��q�;��9����?��"Z<�D����[�h�~��J���ݍD��Au��]�2AÃZ�B�o�7��������c���n{9�l3��937�j��.[�N�_�U��v�?Y.˖>�Q����+��|k�����V��bO����>Qқ;�I|�S�@cS��tq������AS<v]N-�E��+�5��q�<���nq�sDk�4Jg�ц��f^�Y�����`��#|K�K�Yj���\�?5�M����q��+;Y~{�۔��$h���� >����E�9�eK�QI�Y7�.���H�ܓ���}�@��Il��e���hH���2�98-vƴߟ�mc��,��}˥r�O�4���o>��I�э2A�鈅ң�
< �G����k�_�q,������ې�[��7ۯ��u]�~���.A�s_GKW�:�W&їƄ��OZܺ.�Wv�X�~���uߍ�H�����/�Ե$��yI�{���@�����|�5��h�"K��K�E�5���z�����i;�Ӕ���#�q�{G��Y����HR�1�-�
3Q1�kB͏��Ț�2���Ws	��G�o�"R���k��1|��j�P!&��:�l�b�)�����^���［��-�gQ�dx�h���ې�����fb�c6:�.ܵ���,�T��.�y�2��!��A���GC�m����R�l��a��<TS�G
�Ym��[��A������["I�~�i׊!E�|�Ğy���U�.��K�۱�p�I�Z��ol�:�4�+7�r$|E6�����o�*�y�!��'����6������o>�I%[_���rׅ��7�q1|v20g����)���ŷ����D��>b�T[�1ϑ�����m�˸_J��b��9k�n	�&0����g�����J�Y�#����ڃ��;�\�Ol��^�a�*� w-3fi�^�4@�5����:�?�"}����+��h�[�Ը��)�(8�VH�cI�8�εѹ߯M��R��)q�v@,yn��|�@��5�h?g2��8?�}��T��2�tU���n�C��Д�!N�4����y�冥k1@�F�;5�٤ZzfG��wJ��o�Ҵ��
���z�gw�U
��Ql�/�5��[jՎ��(L������ޙ����7����ˠ�v��wA�	����fZI�]]O�M� ��v�ڣ[��"���� ���yJ�����NV�X?��?0<F�@�ko�z[z��|p������=Լ�Ϥ'�N�o���7Bc�:��?N1[�{e��k�t���/�Q9�q���Yg����2̰�$��l��pt����ُ��j��+k��e�z�ϗ'����¤GYj|�x~!fl�#��_�j7=�����O|�.'.|}"jZg	�X�O��%�F*YM��@�"���z:e�<x��!�����OZ�<|�����J\���'�jnnP���(��� ������3�sƹ
p�R6UI̹���+?�\�6�B0�v4���d�䪇���͜��%��z�^����4��`��@���ܩ���1���F�\Ub��D�&�Γ��׏�'�O;��f�'�cn��[�����I9����߉L��P9̩�]W"|��1|�Rt��׷��r���[����k�]�����9��wT��_�Hn�w�XW0(l:^�k"#ׯ^��:������G�b�YZWY�j_Y���$��բl���QV+�T �q��;$/_������;n�
�#�_�Q�dW�.��z�Ɛ�Y�H����<��$��-Ƙ�"�K�Q���B���d��/y��04���ؒ��ez��0������xG<��4�F���hՅ'�[uAb��Y�]n����=�]��s����'ډ�0@�'�		;o��<�v��}ql�ߟL�?�8��yOsE/����wVW�/�Ƣ���
�re����y>Y'S��Gz���x��|�$5z��+Ћa,��-sqھ<^���T�aQ�NlNR��?��p�M�����i���4�JU%C��x2�����}��C�׾`�����D3�3l{� "��Ѻ�Ȣ�U��q�o�Gy�F��'.��'�+
)�D�A���ɧ�׬��b��t�jD�v�	U�*�,��ïyM�B,8��F������ ~���	=бO#�2O1�)�����/�:�6���kà{9ZB�~I1j�<�ȕS����̻[w�U�:!ɬ9����Q9_R;�)rR(`-���0�o�R҅\��P�փc�QQ[ʤ��m�E���w��b~�.`�a�d�Tj[qZ�ڧΒ�>�w&j����L��M�d#K��X̍�M\�{�V½oYSL���5�|j��.JW��ݠ�A�F�^f`�?�1Պ�M�]��X-]t�#���9V3ȋB�@'u�i�]�j����'#S��`�Y��ɩq>t���hn����;��g�W��6>P�ͫ�\�� Da�L��d�

LE��MM'��px��:�ŎP�R�VB�}|f�qk�U#U�K"�O�W�{n��I�>�}�Wmay�/� 
�ଝY�(��y�L�.�R�'���_#�.}�Ѓ¢�]�x�����0d^y�4��������\�����AM�/�ԛ���}�m��X�Y���i�T+���EL����Ҝ|��9g%�n����xh��ݓ�t��}�{��%��67����k��嵋z6x���\���˱��r�{Ue�7�L����*��xZ�>dͻ�ޖ3��P.q��Uԗ�X.�F'%g�8��|VB�ؑ,x���b�k��.��}����3�^�d��Q�b� �.� �EOW��zZ[�����JG�8j&6�5�L�C�iU��k�j�Bo#p�m~K�����!�/�ʑ��a����;�MK�`g�Gi�qX�$���oV�����}�_�>�1�3m~���Q�Q���p�7/�����L�Y�.�.E�B��W	g�W^���o8��2������$�.ȭY�˜W�^Jޠ���K#Sr�$ݵ�vuvd�F��hߕޔ>кnt��p��q����= HKZƟ�v��I���>�f��Ag�-��R:�Fų��&_B?Y��@�O�}'22F��kB�b����<SmT���K��bi��5l����/�W-��ɒ,r�p�'��934%�S��#-�<�Pbg��vLo~�l}���K�M|���Y5�Wg����[ 'ªoD����^�k�!��`Ա�uY��!�S�a�E A����/��ބ�\���C���ѕ�ZU�륻��uU�Ni.��e���گ[mu��gߑk��r�	��Do�dF�5���/Δ}$�T�T*��!}&�q���?;a����)~�k�8���aX�v'��C���6:	1|�˺��~��8�vV9%��I��.��L&�h<��^sĆ9��],�D鿠ڣ��z�xf��� ��;,3s��`V�D��G4/6��n��>cD�s��?u��:I5AR=��_�Kz-Q����B�>H6/,�~ȴ��Bn�/7R�k�K��N_�Y.���φ�"�<eeN���	܀9�:�n��
F�̫�������q���n���i����}�lc����j.�M(x����tP�;}e�e��e�=a@� �q]v�u������.a�i�"��_96�HQ�!�c0�=������˾0��$pMa��[���������?ƄW�~Y�w�=�uߧz1�-q�k����e}����R�Z��-�n�EH����t<i�y���5s�lӑ0H�� �+ ��}��WBDj�'f�˩���0���W�0��f��¸H����%1�_,�'�|?�B4�x3pK��!E��kn�s#��?"����z ��6�l�mX�E�����z�E��>F�����ho,޾���K~���Cs��bff��+��abwZ�����v�����(4ʼ�59t�����Mّ���j������Ldh~wV�P>�|��zJ�F��X�`LX4�������c� �}��8�������0'��+�Ed����I��Qb_��]�D^j>
���f������d����w��M��)b�)2<j�_m>0��h��bZ�^�'�(�lۺ`� (�5�K���d�7IQ�(�ʖַp�Y��)T��e���_�^�3�j�Хuҕ����ݞ֜Y-�Y�qk��k&����LK���o񠘫^U�����Xi4�f<U�ɢJ��=�]Ў���wȪ:C�ߝfy�BY��/T(1L��Gw�#�s��V�Ì���N�kId����_�������s֓���9[x��U�S�?��P�G���0ٕ ����C�$$o��@Yz><U�qa(�gq�	a�J�yg���/X�ś�F���	N1
���D�P��N1���>⡐��[Ϟ6?|��q-��A��c$������sԸy�)�6Xt��s�O�P��kAf����p�� Ѕ1�=����ܱE��MD����O�T�>�M7Js]�Zf�t:����*s�"�s+�]$��+ᛃ�׾�
K4}�����
?������e=�7����\�\fhP��E^k�~��ɋ����U���:��!��T7��ioO+M+�L��K�*s��^�bF\���I�y��TF_l.��V1f�����e97�O�	�m�[��q^01�V�ڴ/�ɴ5_��M����r�3��iU��F���V��Y�`B�S~�z,���p�&�[��و_�70�I���' �gvi���w�O�5�=�>���u;�Z�䷻ц�U�WY��ؗO*����M�>}��e�9�����x�+���
a�d*��G��ƌW��L���O�F��X�
�R������]�>j�Ew�������.�*i	a%��bq��;�0TᩋS(놀)=���iSx�J��v)�4�K���f�<p6-w,u�Eq{V���5D�O�r�k�x��%Z����Ù��ž=��v<o���M��©C��{�#{�b���`/�⍰/��Y� �YIo`(*�K���`��;)~$ϥ,�2��vذf��L[s�ǹ��Q��ڀ�\������>��3����p����?���B�H�F��)�M��7 �rwD}'n} 6�����o��fx!┕�E�n��mj_�*�W<Z�\-����D|�¡��e�j���\�.��>�Ȇ���%���ev�LL<W���b�1|�}�zux�,���c!ۤ����(MͲ�Db�W�OZ?@y�����y����35�նx6A���l��SO3�V�+��!2�a��_C�U@d,'Qy}�l^z~�	�ݫ�`�ѳ *5��eL"[=�����5I��C<I-�ħc�Y��z��SY<��[��!�;��[�?�K�ў���k����ص(ܠ&^��a�D�}�.�)xs&Ct칅ʄl���"֙�'�Ѿ�FJعdAz�Z���V�����<G�Ή2!���0�ｲ����&/Bƾ�\�b�/����6�dC�����_���lk7���>�m�ak�G{tJ��Fwn_s�bܼ.�`b�S�;���q~2���G.2a9>�&�x#����&ƣ�Sȁl4��z2�_麏j	⯎WCI�9�._��I��r =L��En�f�p,;��H	h�����>�zBP���K0PK'��P�Ưt�����^&��h
�S3����S[�Rj/�]��8��F؏7�p�r�����4�IV�Gޅ^������v�r�^��|g~���������NS�G{#��О��)�h���y�v�C��ê:��}��[h�5���G��y�=`�x�J�pv�ژp�N�s�`>S.�l���\�n�nS���Z�Utza2&�7W�}^<g�|����XL��*�-�}9��ȀhX`��y,}d��;����/��]3g�������'S�y�g������>�<u!|�������<����
���qБ�@e$�/n�B.w��~А��u^^^�w}j�[b!����$E�޶�sO�f墩o;n�]��l9��K�J�k)7��B)��� ]�EUӦ����5���>(,�EO8x(,Y�,z]5�x����e{�0�|j��>�'�T��(9缨�R�����~��/��f��Ҽ�Mg-Me�S�l��k�;p#@m�����ZR�R8!�n������>���}x�>�R�1�c+�^�Q�=3q�{���C�H��kR��g�� tK@�L���f����:V+�4��U������D�m��r	k�3��W	���ʎm��-�B���ʴ��|x�|�-�e��7ϑ�.�#.~j7xmo���k�Iw���Е⚇ ����yyƹ��ڭ*O�}Y/J��l��gI�.���/�"���q��i"�Үsg���q�N���V!�f6Ưm&��؉^$�օ7�MRf��$$�@���m���M�O-��Q���r�y��)]F�ׅe���,���
mF�#�7������T_7����I�Vq���Y�fUQ���$3z�!��[]EJ����0&�a�`4�El�*פF�iϚp��1�|V.��,�Z�~��⛴C������P�7��G�������ϣ�u�Ā�F+%)�Z[N~���>DOG`�OƜr�0j��ߓ��'�LNg�����K�g�={�73���� )��[���5>'1��="�> a������_^����D�a��I�BXQ�	U]�P%�Nm祤���$0�Q� �t�%�a�Bz��N4�����ܿ�tK�T^� ��q��Y{��>���g���l�[B؄pvK��7�����o~��E�Y��K�>�6ƣ�|@������O8�H��2��ѽ�:�&�W` ~��O@R�WP��W�o
/�-��`������������vƍ��4��cӻ�'���:�;�0W�g��~��ܾ�U����&���b��+�e�n����[�_���]�2B��W���uX-�uz(���!��I�Zlf����u_'�4�e�ٚ�6�b�%�������t׊c�
��1#� �P$�5�j
��L�e�U��7c�QiUOAj�w��3��x�\-/�f|{M,ǧy�*)�_"�܌��P�e���O�%��.ɶ.���<�T�4B���c#�Aމ����R�&B�p�n����W�_.v�_L��k���R�t�����<��8����(�u���捖��<׎�\y�9)������ʷ� B�Q3�����|�_��8>t�A </.�u���|&�5����*G7&��-��h��Za��J�\@v&��m��6�"F��weNH���Ρ~��4��e_�&���w�������}~�3��=#���ކ'o�z;�R�b'�~p�d�~�&���L�F�[��E�g��M;>��4ɴ�Tng�O��ܛC��n�i�[u١ ە��Px͆�H��k���6���^0��~�O3ӏ��|"Q/�t�� ���,V��%�y�,6�z2p^5���I���5�#O�4���������%g#$Ez�3[������f��m�7�nPj���=���jb��w��Tr�I�ݽ�P����,��ۨ,���C�E|���H��D��kF��[�EB�|�v"�Q�+�6*�-z|�?��O)��2��Yg��Cv�~?>&��Q>)�Խ��N�rӶ�7d>�j��H�f�y�T���ix�ZQ��>Uw������UW&(ǜ��(4��x��nqo�܀Oh�
�@0����Ne���?05)�pҞI^��;y�|t��<�N��Om�.���Dd�9�]���
�}�5�繱?�7&��bBP!AF�Q뻵�ܘ�B>�A"�m�)v�ͨ�-��:X�Z��=���H�QhVo�Ĳ�W/$9�LQA+���	��JeI�N��׏<1�8���l�˞H���#a+�s�i�EI_�/�a_wxl�^4zxz�!ܐx^@�ߥ�U����T*�%�:�{S%8U����	)s���e�������~�� 9������F����Є����jw�FP�)�,�O4�<q�z��.��#��������o����Q�=�P�7;PI��<��uqK˨���Ø&񜉄��с��� ͦb?\)k[o�U�1�y�OI�i6f�|����1����@�mLD�y@������f!ԭ9w	�,�}�B��j����=[���/:97
c��(\������ī�i����3#���୯�?�����]5ᡆ�WV�kP[$pdy"����N����v==Cր�]�٭QMpiL����ha���-�,ZzUE6����0K{N~�F�S\�"n����S���t�%�����A��,[L@Ԗ�ov�-�p"2�S��H�>7y��������QJ.�O��8�ꋇ��6�(�&���;���j��RP��zO2DFB_�w���8ɳa�X�Y�n*唤�c��.����S=�7����^�T��Do�k�����"�S�Ś>#h���Zק>���8�A4]EvWx���Hr0�>A��bᄫ���N���uo���a<��{�?�_(�L��T�;*]��I��/���J�M�JO6x��e���11<���"q�'�}4����ͻ�;�M���$q�8�6������Z��R�L��#�hኩ�GyZ%����w��3���_�w����Ǩ��_K��y+ �Ә���~��z��7�U��5 ���G�M���U�D_��~�Gak{Ä	&�Z:<��	A�R���'�?�I�7ij�(�|��)�D�6˸Dw,�ʹ�I��6߃܍�f�M�Ԯ_���}C���8],Z5r�^'�̒����$��	�e�-b1���������H1���υAc�l�BW	5��v��z��*�2�F/���ư��H[�����9t'�/�8���u��.1��Y\FH�;��Ct��g�l�D�ϴE��;y�<k#ˠU�������};ɰ)Pܷ+#3��8��zvQ��oT�$q3�{��Ω�C��g�(8�0f陌d-Xfj� H͸5�W˭���v\�}����a��O� l��6m@��O��/�"�6�_K��w���ơ�v�{[̕R��d�X��ݏ�$��VT�jS�Ϧ�Xɨ�+Kg��������,�>���lc��]�~�Dnf^�9g�@(e1t���-�{���#Y�����3��3vƧ�.���9�'��Z�:�M�H%��(�vJu���ʯ�,��_��]bU
��׍������uk�$z��c� ���S����g�4�;c��Gow(�	�j�@峺ؓ&�2Y���U���m��;����Zkc��Ԅ6F��Ww%����]:ݼEo�mJ���h�=�/�֨�ʻ�~w�㰞�ڣ����Bw ��C��Ǧ���y��	�z`��V��w���(u-�Boy���E�i�̓��s{�;�Ñw��Y����mh(uQ�������e�P޲��ğb�C�i[�]���K�2ӄ I���Q� ^� ,_���QU^����S��B�^���3��^M�ˎ��Ro���2�������d�����ZmU��բ5�Z���ڵkV�Z	� FUQ�R����N"�S�V+Hb�"����_�����r���{�s��s�+Dq�<�]��&=���ˤͻ+&O�u�fߎ��t��<~Z�l2J�<��Ws���_j/$!��G���ޏ�$;�z2�C)�>%�C��O6�Ylwwl�����E���z�N�1V�[E̞�iYi�]`�IИh��f�������/)��%�=뺨r��(�=��ؾm�_ڨc>@etz�y*<B�&A$�=�h;�P{G)�d]�����3\}Z�P�}4��)U �^��+G/{���c�[�6-���c����k�����霼���\FZE(�⏍�Y�QZ[�. �H�k<�W�͸�]IS�!"W�R��uq�����9:�P$�e~��|9)Ǐ4��\C�"6�vI�u��|���p=[���p	(CN����"�v�Q�T�T)�����|�#����F> ʙB
\���tfI����ޟ;�T~�z�)�������lݏeA �/�ڵ�Il��p�RP�[��N~n�U��=u|c�+��M���*��`+���%3�U��`���!��3и����'�%����<m�X��L��YZ�\ ���ʇ��5���9A�9���#���`�Ѹ=��E���@v�KЈO�H(i[j���=�8�3w�h��R�����t�H2����gh���GN�d�y>݀cD\��߬�������M~�Ï��	�e3�	MQ#� �I�2�<�(��1 �n�rUsW��^�4�/�rh�2�v�$"^I��,�Q���މ��؎]�I5���O��D��w�����9�$d�̎Ӱ�DX`>���u��XŖ�˲�
�]~�d� {�t�N������n�����v?�`���N{㟿2]��[�u����n�C�E8�NA�p��јO��kևujq�����w�H�b4ؾ2Ρ:8�n�p�۬2����A��ߪ����,���~���;�f]�{{��؅Q��ѠK_>۰����U^`����6z4����/�<��r�Ń���ScSk�G�Mv�ɣp���KW�~�_ȿHzx��,
�JH�A�@����5�S��$\�rUW�J��X����[%�e���p������".@��}0mh�q��'�WNo�el�r6�Ut)�l�|7�Q�Qy>U��:U�P;�����Y�_U)�$v��*���+��� �@�� b}"�Z�T6�?z�;0w�LS [��?U�f���X	�y������q%�"�_�����jQ��W	m�kk�P'�:��=��eg[������5��%���]~˽��QF0��[���gE+�?�΅9B��C��3|�J�-�J{r�=1�b/ǜF��K2'zl��g�[�����zU�������x��NX	���O�;Q����/��F�U����{|��j�X8�kq�P3��bq���RY�h��i�Y��;H�;�)�f��j�ɒ</��=�Ĳ%�j|��$<p�p�� �o?��T�~'�Þ2^��l��@�@f_����Lץx���l
Ʋ���7��+���1=��]<��TX��q��ĵ�7�߷/uc*�[27�8��{�;���S�B\
d_�_�\�<��=mXk�1=7FV��즒O���L�2��[y.p��=ގN�ܕͿP 7�M���
�Vlie�D�2�W,�V�m� ��TrBŦ��N���S�'ܲ/@�z{B����-��П�+�H;�c�eG�����bf�%T�����t~zwӰѢ���Nf��wㄗ��v����|V�x��[�a@CXIOT��~�K;���;��ˤ��4.r	�+:Z![}I�����']�&�}7�k}�I�3�K���B9����]����+v�
^�K���,�M�jR��/���
��/��4b�����D��Ѵ��~���?�K�$Ī����A�V=��cb�ۧ���\l!pd����L��48��~X�"�>��a%���n�+�c*x�r�>������*���߅>�c�8�6k93ih��V�e{r�^�W�Ґ�*m��[�?Mr�����i�K���K}</��1z�}��}뼬���];�u$����W K�ru3�������b�cs݊�)7kP��*�e� ����!d��0��M�����+�wD�B��E����R�:�a��n�a���<��)Fլ����!Ƕ�R�zL���ɀN�@w���d-��1Á�uM6\o�,Lվ ß;=�����I~��˻n���K>3��G%�z&w��߼���Op�nO>�8}%��+j��W���t�ZSo����+����"�#�o������_�Oʼ�T�����sv/�
��0�M:���v59;d�R` ,]����}�A0��V6t?g�H��.?
b�^!�z�t'�n�����xt1*�@�l���Բ�����Ti���ۣF�7��%����2ʿu�β#��.zgO|qw*�3	���pX��w�ع�|.��|�{�ԗ|�����]A�L!�
�7%j{(rTh>1t��[�)�t��C� �����g��U�1+hw~�:m�� isb�]��z����������9Vwn_i˯<����4��I�%D���`�&�������S�UgoR ����>�_#>vr/6���\x1�yh4�_��5հ�]��0.�#�����_׉�H���mۗ���6�	̇���&{@��Q�O$]��z�Uh�|�Kt����[֭�j�UO:�-���C�e�d����'��6n���Y9�������+T!�o���h�����)ִ�y��/ar�hT�tFf��'M����.n"Zu����������j�����1%��0n(�KE����[��ш:/���Z�5�Z��B����J	r;�~����V1wZ�?��!����!��3s��z�l^��YA���K|P��:O��j=��Տ,YF�ypr�(6�b;�z��Hw�5�.�|�'hR�Z0$!�ʣ�{�~����~M�N��2WY��ڸN�d�T�Y�GN�Z6���Nu�����ˎ�ɲ��W�T�p#���9=�ڤkH	�p���nu�WRr�QS���w��b��5��@=`�_�DFF��?s��=�4:���F�8�A!�e�߹���o*�
���\�h,�&��q��"&$��Ȩ&�jW����"�r�f"����ME����o�VT7M�6X.�ny5?��/��M��)E)��
���0��?V��}M�>�ۼ6b�v;�8I̙%���[�U�s4Ռ��7Ҕ��F��|�n�UF�]E ��]���鍥1��ӄ���(O�����鲵�����y�G�P�%�r���2�Sӧ��ɝ{ʾc�>(���� l&`�̥3&˗��#t����nH+���ef�"̣�؇%�c�ء�=Q����}i^���~��n�b�ڿ�>ק&�C��biP��ָc����a�ޞ�;&���Xp�I���^t�n��S
Jb(l<OE�^�_m�_&e��5p����Q��\��L���c��gָ��i7u'-�$��Ն�"/�W�6d��!Z�D"��Շ��?��4��f�>��,�f^ �H��T��������٨���w�M��e��x�I�<W��n�h���#�tMm�9�}�5�K3k��6����2c���q�*e/8���h��^�(�|C[V�)W<�����f%QK|�Q2(�^��d.k�ػ�MIf�:�Nn�;T1�O\*�����B���v��,Q[�@�}e�Ax�>�=�t��cV�x��R�D������=�W�������`=� �!�܍8�'�@l�D2�J:���Վ+���G�؞G���R�-�g�R�8�o'��V�Rt��Ͻ��Q�H�UޕCU�P �^�v�$-�;�:��&;��=|�D^�8� -F�����n9�W�(POd��udy��N���l�w�`���/p����̸P�\�8��a������2�W�8������{6�~��(� ��\�L_~ҡd�5|@*�	�*b����ԯޫv�۰�ꮗ������0N�p:HͤWI8�� ڥp�Y�Yn#��i0l�
�l��{�WN�l���.��/sl�{_V'}��3#�+%�NT� ���R���Ŕ�$��%h�V��&��@�4_|��~w3A�K�`0~:�;1�wd��d�9n�1Ujy����W�T����*�_���t���	���%ձ0�9����_��u�݇��ۧV�PW��&7���'���}���7�R�n��N�)���Qd��s�;��?��w0�ܳ9�k�*�QEX�����.X\�'�H��[��č�'�K>l["�z
�����L�E3�=�+:�"��
�N5�Jӣ�̤jS�X��z�fvjE��_t����9�m!�^�\����d���A !CmygO?���v��	����b_RY@�&@��mng5��^�ۺ� 	��=�#F^�̚!J"lo�yp�Қ^�� �n�9:/���췦#0��}�_C(l49�7z4�7k���SGG 7�Df�I)���A����M�����"�;S��S�O���Q֖л�l:�����PL
�}|��DUs?�����uy�OeD/��kOf�ˬ�r-����F�6ۘ1]&�z���e<��{Օ&������ܪ�[�+5K�}>�c*@�I\�Ito���<K����^��_p-.�~�"m�t���Ö�a�s5u��j�6R#�u� �5��:ӳFWA^��~slZ�{'%��x�D4�����4o�׏�7�ґ,�Yd�̥� �|?˪omؑ�x�+u>�%}`4�����6*�E=�~�F����r���r{>�O�ɸ��p�/S�M
ݰ��"�V�&���e�h�XH��$�CJp�3��@�	�ec����_���`�'�a��9�'��~ߩ �(���.w�W��+�\�
�a����N��mU�xד��U�`|�2���&�u	�G?,���Wԅ'4lz���4.��V!�������UA
נ���U�f�BzL�4����������=E��޳]R2�!T�mk(,�Y�y� ��4_�������u@D!�4�"~,T�x���@�a�R�<I �����kZQB=��LG�T@�dڼ��M����y�
�UNT~�@r��˥�W�z��嗣`HrK_~�!�<�UpZm�]���0�(�5_��dD0j��f��qeO�Wq�S�-cZ�������2S=J[H5I�wg�{����݇�t4��_��'��F�C����q���{��!��78.����QlJ��I���O�Q>7��3I-8��6�+\�0X�ީ� 7�����.�⥺�N����Թ��� ��F�g���S[xq��;��3]��`����8_��� ��Ȧ�
�kΡk�K^�|�TNQ#i��]f�7��hh��Y��;�>��X�sC��7�~��:����㡼wt�.w�G=6���δ����̶�'v|q<�������)4�)�1&sU>��V6��;��z�;���ut�`fSBF]+��ⴀ��>,ό�)�r|-q[��ӗ���
d�Z/��5X����*���1ZΠV��f��5�R�*�f�MS*�˱չضQ2��@~��=�[��nv��܆�b��n��<�/���9Gq0�+1�n�X��aAh,�ڄ?C��v�)��N4{�e��?�Q�[��+��n��D�v����k�?k~ࠎ��2�=��A�w@Ew ������<��J��o�ןQ�]�7dg-^o�t}]&���������+R�󩕖
�yk�y����4=!<��ia�F�1���n�i]��a� ���7L�)�Y�b�V��n5�D���w74O�7�y�m�D��ˇu��/���?Ny(�����V�m��Q]�U�i��߹Q�?���|)i�-G�1�"�*�žSux���Ygab�[��]�	��@����c)\F��u�'z�Rq~O���4��Z��r����t2]�dI���f�'�����Y�_Rc��qߤ��,�w�1Ήk;k�3�"���J]�WOM�\\����FNߛxk3��;f�ϊ��Y����D��Ԕ���Z��PklOw��[��c��P�ά4�+�F�=�R���F[@�����\[�?k1AD���4عh#a�|�K!K>4��5ZT>.�\l���8�a?�`H6�NA�1�����P�����	Hsn����i�L.�W��9���	i$O�5C,i�'=Uf��ަ��p�x��\GW��l�q8����u����/B;�Ӭ�Y��	�6�0ЀY	�H���������1��e,�KNs��lw���X`r��ՅH�6鈆�n�Uf�A}��$7@���O\:z��+<0H�+]��J�h��U�"�ɶ�� �����9G�yF������90U��!���<I���\z@>������ ��;cZxN���,2o5aJN�p�yp5s}ǉ:���MA��:�C�eb\�
~�&h(%-��e-�"R
il���ղ� |a���|�G�tw�<�1����@�r�}�$�Oԃ�[̰��Wi63! �-�6�<����#��:�%��a5r.�9����R�hn4^O޺8E;��R�%�Q2_�ҧ�����_$�$(Gq�p�'C�ni�wO�2Ms]�ΈK2}�o'�_�����@�k�G~�W>��c�s�7�K���� d;���w�s4쫵v�b�b�4�,C����0����P}�*@f\��vUO����^�Mَ�hpy���[vwm�ӫ�X+$��'9n��a�c���u���D6D;o�~�"Ky5�;�#���n�D1��|q���C�?�N˦�6������I*՝��7{��������:Q2�^;���SB֪H��(ݞ���|(��y6aa:�����`sO\
����K�� ��o�Xz�Y{��O�or3����|}��Z!�����?Gz4�V �V��c�O.�ȥVcll\�шa�j�7'������|<�W�Ƅ���O�J��L��;���>x����4Oo���*�Wt�Ҏ��?Kڢ���D�&rS����iņ�:��H��	i�O�)U8��\�6����������[�Z��tڜ[J"��vjE5����iMf���XJ�{�����TT����l(���b\�"4^f�a<�n�S�òXA�6W�����u(����=(7Q�z�̋�<C�dU~)�/�e}�_'ц�=cxE��3�&IPh�R�_Yi�}��Ӥ@����+Ѹ-��E�DtrV�"�bA�(c�M
��iu�oP��Y�zE�#�I�?ɧ臺���EYM��ǏP�kS^%w[E'���h͖t���2�>���Q�F�χ�r��I�'�J	z�(���ׇS=(�m֗�IPw˺�ݘ�O�e�!ɫ Al�I���v��N�s�`0�<�@�u�e��1��}�gyr�w@:��Q��3pe���^{�Z�9���������-���P;��pL����NƎj���wN!9��w�#(lɌu>o�>,L�G�����_H&�����������R�߮�1ߨ
I���f���D}=��n�V&�#��c��n�9�"K�(����b� $�`z�b���կVf9�tr����;ƒ����LM����GP.U�=7�$Z�WWv�F�т��L�d~�hn��7�l��%��w,���u�%�����'����lX!�#_s���nn�EB�mxngHlu+ڔKu�\,yN7��BH7�E��S��4���<Wʲ[+l(����.i���gڭ�� ��&�}��Գ�Sudb��ͽ8[�r" H]5�h�=�$ lXߑ�N����'ms����¶O p�| c���h5~Rv� V-G_�9J���/��Tђ�6wo�u�vn�3���(� ����k���ad����}6��*.�-��-���?�/Q�1��(�Ŵ�=�طH��,�1�~k�����J�Y� F�M��L[a��+-|�+g	��X������k%��5��Յۮ��{�)~?6�����Yk��9?�B����{4h�q�Ğ���������`B�rO�(Їn�@Η�d'��x����b�D����*0j�yy��ԣ���[S�k(�ڪ�_�
R�r�蕣q=~Z��r-�ͣ�rZ�����8C,��׾�����Tk��
��w�|�	!��T����Y�(�c�fH��ʕ�8r����K��5{U��(�m��w�3B L�pkm���妶�Q�ۮ$��i=�n6��CP����:4�F�U�����CCm�ʨ6���;m!�6c�=��v�b�-���_ݟ7d���'M'�6�U��ԙ$��f#j3�:7�H�7�v�2��=��?ޤ{N/j���xk���0K��������,d@��sbh��F>�����n����ʢK�\������77�{B�J�/����_�%�����Aa �ғ|�S�$��E��vH�
�.Ǟ୅#27'E���ބ�����27�)Z���&�@��d��`8�e8�'��x�5z�n�JX`��S�b�-���VXt 3r�5�"���p�"&2�~��E�d�<�^~�9��kv��f�23�m2\�:�%�~୅�� ��$���qO�}�jK6!�.0�(ό4��Mr(��A� ������&��`���`�ds;!*��eM[�5�,8�7�_j�Z;g��ܜ��f���"���@s��<|�����%;�0-�k�mY�P�4.Px�+��1(��FyE[���ԉ7�f��ѫ �_짱���sn;q�/k���y�	�#�h�z���uIQ��D�]�ji/�"Ѹ�xT{�[f%2d�6+�Z%zs�퍑ai�HI��*��2Y��}�n�^T��A�#nRm.��0yV� ���X��p�X?���:Y�*�8�/$�;}i[�$��}i�O��G��.q̀E?!��v������X�q�%���/<!�����yAĢז���=Fy��ڏ9 @��F9�jF��'�(���ԁ����{\5^t���E�刄�opk��Yz��;GEir�m�I	�<M�K��7P���1�T}�{��%��p�䭻Cw�;�?���劸vw��'���X��ۿ,��1�"�o�ǋ��l=��r�,�?�Mǉ_��Exĝ�+K���; N%kf�{���[E��t�b|���B��2���	BA)lza ��w`�����<�����X������v8��i��A���;�4��/3�
l��Lz36|#C:*�xIJ�,$�����c�H/A(x<�`��\j���b���󚜱,�6i?Z���Wq^��c�I�5E�̐�E�Y�U��Wvz�b'	{<��y��UKO;�%��]iH���slR�N���jY}�
��[Qhqz���p��E"�����CRkKw��\C�)K`�2��n����/S=����x���Hi0,�����N�����/�<�P�ke� �2���^K�-2n�	��SLg���sWfJ ��G���CA�+�x�A�0��pqu�U��^�P"��f��j��LK�r�'2��1���F����5� k��Ý
a4�5u�$�Z���'Ĺ|��^4�a��!S���I������ꅗ�xV�kz仝H	�8�7E��g�/WV�ퟒ��ў�̗���"@Tm/C>�-c��~H�;��
=��"q��so��P�-�+}L�r� W*��A�����g�{M�A8|`�b]���A��R�,=�|��6w�����_�.A#Xؠ�_T����YHQlD���j�h|�ty����x�mZ�D�W���'��S��C>O��&��"�#��҃۞$5��&�?��l`A5�g�7pm)�ό���6y���]�fN�#T�1p�%3�(,9����zp���Ox���>gRxX��x��06�T����s���w�s-�UF��a0�y���&�vbD�u\�?��`�#uB�iCQ��8.%I\�jS�}E�����z;[ž��%�w-��xa;k�!\�TJ`��$3NbJVN�WZ� <B ]`/����AI���>�^x矾-�z�T�?5�{�<>;��k x���e�����AĨ��*)�s^C��10mP����������%�U�_�ݽ��x�N�_�Ұ_1��G���`�����@���O�I��&��͊��+� �,�VR_y���
2��R���h�j�.c�a�b���7l?��ʗ5��R~;��]�wz^���G��L~Bv�f{g	e����w�����*���2E|��S�dR�18��(��=��n���L6BQf�R�TJ�>�`�M�i����|��!	�P���/�0�B\C�B+-jӌ#�G�`��r9�J]�p�ڞ����[-'M=�"���#̸��U=!x����9�ap�x�������J9�@=��b�+fd����#"�z��̙����2�gD�5f�\�}צv��X�����U;UF���.�07��Wί,���<[]'4���yT\$y�r�G1���h!a�ݝ�?�>���7ގ��1?D��Xj�QS�I��/혚��i�����8�|��L>���-��t�Q�r-��}��qXCQ�ˋ( O�Z5nb��狠��;��O�X�f������tS�y��V���"�������pH�~Wm� ~.�c(��- �ȯHa:�����f��fÆ�J,֭�ԯ<�I�eε��sۼ*�e�k&��d�ں�B��'d�Y����"!+dy\疃6#u��
��5���L��#�Z���A�L��+����v�,�8�]�3�,z-��|]�OF�i(B�u)b��tu}��O7�u��؇� ֬�#��]o� 3�%��;�@̄ol4/.���G5���(7��4mc��HW�FI�8K��=���_#͞���E�]׎!�)��,ZJTZKT��Ϻ�>���Ce*~�fQ�2m��/u2m���aԉ�}w�H������AR�>��M���� �iL�*�iWS��>Ų�{��|
r�������������Du �7[Ļ�Ŀ7"@��,�|�i�9��u���� 
7p]�̫0��B.i�z��[��ޱ���Yկ����0��D�>?����]��*��#�p:x�WUS}��|V!��N��8�l\�q���&�$i���c������-��}�"��P�_��g+D���Vw���^Lj�s��,FM�_�F�<����'��7H��M}j|�K3�����DI�[���eї��oc�;=��#B��yj�1�hW �<�4�c)`	�Ӹ﬽���ܖS��ӷ/=�_�*A���th�"/���_)kn@]���Ρ�j�� ޢv������{<��+��9�??P�=8���8�~y����VG���n�^ش]����7���qw�6|'�f���H	�7v�fl�m����1��+�ƴ��%�\(G�d[@�_�7]$I���Iй��$�*�?7��?)d�K��������(&&���+���q���r�`9�M��0�geHԿ��H���98�(q�ةX���Nۛ��p�c-m�	�aE�m����%L��7��j���g�J�H?�,;�1�DѻU~}׏��f�RQb.� ���|���u��o�n�����3�a�"OO���j7����%����c�ҧ����-p�今^|�N�������2���r�4�3��{��׎<<��=��o:bŞ�׊�*�~��p�)�K�~�It�W�D��;�l{�!��=��i3��Y�p���E(�	�U�Ӈ$FM�ۮ�F�q<�`	-`9��u��{"��a��m<l!����;+)�:�QIDCL�#�D뷳O���UŞ�W�n<7rO8�c�
�}eߟ���1(��ښ{�i�����.�_���p��%-Ѷ���s��Ie�D:Ŏ����++�y�9]��W� SQ��~M"I�>��Ŀ�8�Z�I�AW����>��ܦ;�)TW1XE�Hl�X{vtd56إlo4�V���/Gܞ��6�&9��yӴ�g>��r�+�b.h�$��t�/�ݥ}i�
F��9�?�G�##-}���5C�E�Îvb�t-�N���/џ�|��ʑ�:�)RL�1xzkT��ĝơ%0']H~��v ����_�ؿr͂D�U1��D�S?�`�t�9��t�cK�N a������ �N�"�Q^�3����|�g�ԇh�}n�y�ˑ1V������ٜ�d�q��V,.C�lt�4@�������;b��oSi?�8��\��Άx��-_@>5K���U���f��v�����MW�D�� ����Ӎ�hz�x>'+�%Jm�su*~h.aG����2������_����0�=s�>8!9^|D� �V�6����l|�9c��+_�}�a���Tͫ����&��֑���ˌާ��w�Mz���j!r���"�3]�[>&�?^�ʧ��hن�pY�ͯË�=5`��$���K(��!�WH���9�OT�t��ь�*O"�f�`7��;�;�T�#N����T� ^�{j�?���%�hX<��;�%{���A��:�Tmk ߴw��^��e� >�?��&;g��� ���U
\��P�C�!�:��c����5�P�8��cڲ����h�Ӈ�`+��y���]W";��n�����Ԙ�F�����J�PY�
��|vvg���b"/N�ӧ�B�k�����2	ߨ7O����>�N�7��W�tnQ#���p��:��C��Q��Ϣ�Nw�C��X�'�ֵ�\d�Y�{�$�w���}*c���_m�N̓�"0~��1�sX�Q�^$f��L���\��dk��Q�<������$gd����޳���I�]}�=��S���f���k;��5����"c([2���y��"ޘe[Ti�n ǚ<�ä�����ݟ-u�Z'����ٝ�Χ���*ߖ��,T����Ut��w�v�9�-�w��z^�2-��g3�;�c>�ߛ[$�-��Κ.�tۮ0^��^=O2L�Ů۹Л���A�d.:i����[@�����L=�8��Y����1 �Z�X�8�M���F�����E�rRa$�k��r�;/@�C�&���>,W[���i�l��e�=��?�b��(��Ұn6��-5B"��\0���e�z�L, ���A���|8��y|�:�G�E�Kn^x�U�(��5�d�Z��C���ߋ������6�1����������.W�0�d2[��<�E`���Hn�y`~����yBvw'��P
&mwP^�3T2d�w.���Y��f��zE�E�r��yf#	��.�A|�SG�\������n=�C'�m�ç��+��>��25�����'v��������z"�i2���b.X83`�����v�nKFd>�9�X�%^�Q2� �ᷗǯ�
�{-f� dԯ�X�sKv�G^&�6�����2!�U!�3(��A��Y���g!!O�΂b��qeqK��?��1�2?�-ɢM��1kKc���r����8Il��N�A��_��<�w�L��Z�΍)��M��VߤEw�#x�ou��[b���#���h��?����76/`�g.�Qo�k��"���������g:Gbko��}Њ�y��3v�6�g�5�iwC�ycu��ĵ�ya�_N	�%�nX��U��Ix�Ѥ���c�K��HLA�1m�4���Dl=��i�Z��S��yq���[xa!��h�&~�����&07���g�;�eL�7$AFt����w�Tp�6�S����x�7`W,hk��P�P6d�eg�c�wƜX����{�������j��#�g�.�N*��y�#�_�r8�� Ҳkq������y~��jcWu������B��[�R����wty�`���!K\�
��`UNo���{�,А"'�o�]/_C���
����lR�U}d?�;�?���941�G(\���4|�������n�B���g��y;�Lrٌek��e7�Jts'�9ρ�a��>K 
ʙ���L�M�m���Wz����~yO�� ���31f� .��yg���	��HO��s�Y	�U��x�_E���7Q*���ݪ�66��{Hd]����_PI�*y�%L�r'���8.S��AYa��䣩޾�7��� C��"���M�����I�濸����3�v�C5��(g�Q�����4��gȕ�����������`&��VZ��r��'P��ښN>c	e���Ƶ�188K�����=�(Z� c����3eA���g���w&�|�50���Y� %h.14��F���~?�TM�x��{�ݳ�&��v���@ؐic2��Co��4-@k�y2m�77�IJ�hm�0c�Z綖�xB �xB(�;<��6ٚ\���
�K�B��fq�N̩���"��f�ij��;n!��
�y�d��W�ɸ�&����$c�)~�5�\lS��9��~��k�;#Ա��!p�,�ߗ?��}wBy5�`nā���
���"�V4:��E�kZЉ$����H���ѭC������ɹ;�Te�4/C��;ML�T]�����q�1f�'�omP�=�%X\Y�n��C��cV�!�Y���8qG���@:�,�,)4�\i�2�~��0|�~z�B�3�=maX��^�R؏1�I�����1,�-�Y`�e�;�-K��6��,�4у�̸_��ְ\H�����73�wj�b6�t.Qx�v��1���|{�K�m5�q4p�~HH��歋�0D�'�z0�����s�]h�Ȓ���E�� ��:(�ܧ4��]�,���J�)�d����<�AQ�j|�0���VJ�=duX�����I�}xI(x���`?8+,�s��*�?#�q��G�:�dwԻc:R a�K6���zy�D���9;����^0�3���,�����W�������{u� ��/n��.3aO�\�"R�R������*�����;jj��q�����z�'���~�Zn9Yg�`by���H�ױ���H��^�1����q���3�tyt���ܤpz�$��GI���殧;b��y�^5>�h�+P#b<cW�?h�?ք0~ 7�i!?��s��h+_fNw��H�4�r�j���qAD�/�O][W����F�����+~�tYp�9�xp��׶H�|=M����tQ����JMAF\[�K�\����%�(2�Q=��jm�8�e	��T�Q�έr�7�w�4�,#��c�J>4�*�'M
_����h��+�j|^}3E����­Ք�2j���Qk�W�9RJvz�y1�v*�	�`��{�#����s�Z��d�Ə�l�����-�²�q��ۭ>�$K�����&/s~��ϸ-�T7��a�"��rU��G�o�����_#H��1�/6}�vA��w�/ߞ9��ví�n|�%v�Dp�OO�XͲf�s�f�@�@�x�n�Y ��3Άo.I�q�%?s��U�=V��пw��5��V�,�]�q��VK�I�0t� �N��TԼj#�z��ۛg��$
h�4
 .>��V��glt��K`EMj��'��W{� �%��x�� ��R��r��13Jv�+�z�fe"���G>qy�?�T���4���X/�.+��ױl��*���h@�_�=������x]�R�P���cTs1�F�ɲ�k�z.@�B���`9:3���
#��u�[c�l!k�}��ZJ�6����!pC�c����7��EQCdX��lj[6�K������lY<��9'���fV>�i���o�)G��D�5�C;�o�����G��>^$�i�����Ûy��?mB��%�7��eh�|�Go�TI,��׫óc 0�f��������Y������=�&3�YF��D,dQ�W����n�U{W`<����CT>��R��)&/�ۤ-�t�h��]V�g㊍0���vg�x���H�I��W�_�aH(`?}+�g�ӥ�{qj�<EE�D��Z�e��goٺ[ş�a&Ӕ��,e�۞>�;�Q+/�Ν�U�G��ܲ5#�����M��e ��������n*mgؠ�T39�%�C� ���> u��N���N���x��Bp�q/4�ú{�����P|�M��b����yr�����v>r�j���^�t��*Y,�u�d$�a(A�Z�X9�s�<Xt8F�������<���(,pH�k�z<���L=�e1z�HVa�$'(�Y�N]�5��@4������ˤI�rX�:�w$.72$�-4�h|�s�Tk�N=�wOL;h��N�&��N�=\\�,���:Y6�j���ɥBY���ٺ� �׿}\�Wi��%Ϩi�i�*ü��'�ú�k�ǌ��mT�B�/�I�1�ύ5���=�7Pw�v��'���֮�w�Yp��8�3K���9V�Km�S7q�A-�+c���)R�����dٵ��g��Vg�8��q/@Փ�ZE��2Τm��ٔ��X}�kL�a_��i,���o��B�md?ѣl%�j	�� C~o@N��P�Nj�k��gn��������a7�[p>�\ �d��X��`u�,�����f���J��O�6��s5��s#��h����:���x����7��.�0>
����z���]���D��u/�]D��䓲��v�c� �����>g�'.������_מ�:���}�'z�ω���$�M�����T�d�=�'j�q'�:�?���|Y��,�*;l�}M�V1�@���`�e��2�+�"+L[OO�����~��8b�� �U��������J�:B��B�!�J9�"1�!1g��9���C�P9��36�D�q�4��|�m�3~���|���}_�u=�}?���:���r.��h�H���u�?([��:�i|皚_��̙�5Jo�,V]�O�Ԟ���G5P����,����q�V�����������=!��N~��L�O�ǖh8J��n��)��_O�~ù3�!JГ�wy�v��ST�mͳ*�S�̀�:��3*F�G��E�D�)�Dw���N��]�|�����̯w,fqQ��mw��
�Z&��sw������>G������n���^����*C��b0?��S�x(K�tZ*y(�X�ɍ�'�vKN�t=�N����|ju�4�v�J�׼�]��Y��_2�)>}�u�칦��̪Cq^Ý�5]����~&� �nz궤��Դ0�p#��ZѮ�6\�OOĞxv��Z�q�z��%��K��t�28Xt�W�pJ��锳簿�����R�/�Tl�:��s��|�n�~�[�-����[�ŝD��~0������l���w�; B��j�g-iA\>[�z�H����|G �5��q��^6�ƛq��q�)$2��5�r+KG��c�+*Ed�2=��fI^����~��%8�RR�/!��xb;���0���V5~p|�^��,���89	�����]�p�Oy�lפ7����@���8 ��cf^N��oYI\���4��tkޡ�w/�
گ��S�>}��Yġ�j�����K�g��/�gx�uD>0G���Jͷ�WF�2*��"M���B����v�L,���bs�)��?F�ڭ�kf����yH�����L7���C���R_�yg����?���TJ��&i��Z�|D�|��E���:��Hv�¤��0�v_��|�N�^ԩKTQ���%OK�H�x��$���[SUx"�zZ�ܿ�N
竒�u���0��| ��9t#�����2D��YMl\�"&#\��/v�ԕ�3w>�x��.����ԍD����.����w3R[�,i�CjW� ��[yT��jD�,[�H����;d�EPc�L7�ז0�
�Vdl�s �K3�.�dձDX���X?�H�]�N�,t�Cd�[�����"���W�;P��/��(��.�Q՘�ؖ ����*������w�*�^���}��hޅ��>���G���w�C����]4���+kz	��R�pvn�9��XH��~�\zwSC��pT�ş8S;$�V��zc�@t������?8���{�4�v2c�[.V�aI0��\h��~l�DDخ�T�%1��ދ�&�Ş�v3j�JJ�R�<v�;�׏�)7؁\�1O\sa��T������_�:�U(@��<+�,j����sȌ��/L+]�sxO]T`
���P�:�����;�7(�p���X�fI�Ox੠��fs�CTpz�j8uE�]��(��)�9�P�rlzИ*�ܪ4
TИ�}�˨������*$A>�@eˮӡ��ڝ��_�?���ԥ#V,�ވCLZ�$'�#�r��u��1�DJ���T��m�e�8_8��;粞{�0&����{�m�Gӭ�ouVv�OR�����2YUN
�Q��0Y�Ip�B9���I�D�>�>�S_y��xܿ��$HqӚF��!��2��W,5m�G��,hWk��`�+K����f���)�p�y]����QZx;�����w)��)�}Bs�5 ��|�2��V���< �����"_έ�����ⷔ�ďE�=��>}5��%;͗�����K{����/��Z�����z'
���]jǠ���T������O��t_*;]Ӌs�+��Y����N
��!@u�%*p�{��	(?dh
+�G���i�I���'6�ey��,�/���/�����Pp4wƾ�8-�����
I��S����i_�KQD[Y���V�������'�L���;��dq�㵋M~yXiz�0v_���|���a�[);,�Q�9�7ȣx�Uf�ԛ.�3>�W-�U�w�<.܁�*�Q~�?���#+U��� bm}����h'4Ya��es�5*1�!"�ϗ�&&��x��������;�dg�%��!l����.6�����<k����!�^y=����u�Z��Ɨ�����[�]z�?����v^:Up����{��$�5���?�Yǲ�:6<Z�#M���!��o�_іbz��9����d��.�x��kZE:��9"�A�r>��[�2�E/D��Fe�}�st"�Ъ�x������f�/E������a
��)첀=���#�T���c��h��f���j���!A>��� �EP�`k� q�6|8%�wc�t��w���;��Т�Kj#��ճ�7�j��1-��8�jm
Ms����%Rx�����ݼm��{�����o[;���/R��	��+3�}�^����eR�]��tZ���Հ� W���~� ]�F�c������X�������SO�"��Se����C�^	7��W�Ao�_x����N��d��<����p����(!Z$"[��q_J6�/��[P�<q)|����[)���>�&+��C��~)�`���Oz��HC#/��	�s�;�Y�q��3�q���#��d�ߣ����u� ?�=��.��2T���"eq?��@��U8�S�q	�xT��`�ZƖK�YO�Q=G�a�^�[O����=J:�tZ&N��{}|)H$Be�0x��Y���5�$��+��P4�ks� ���2i��n�������@Ϣ����I�}����b�X�B�`>_>�4�3�[��\�q��j �GG���:�󟈔bL��$�~��]��7L�Z߻d��y�j��UR�J>��ּ���4������4b{*��EB�E����&rR���9����u��w��Υ�U
�u��^k*�*U�t��:��C�d�%w��ݫ-�N5��O)�����\��W���2�݌!9U
#}�nM�W�#~���j~�ųKѐ.�nr2j�h�A�F�0��&���w2���o����x������3
�]~(�0/:+1��l�?)L�I��'�h��渆����0�)��#�KT�uh��^�;d{b�Y��$�dg1/�ϰ]�[�xU��NV �|Jk=Uч�q}�a@����$cKh%�Mt�[��駁��<����T��CM�x#ޟH�U�n���A�G=a�9���+�l�<Z�ٹ��4D��{J�*N0`��'��мٴ)^�Ϣ)���;��%gl�We���Q+�
w&�w|i�'���A!)��XZ��A�E��k����� �RaN����J�4�9JV�Mú��)D������i;�|����g8֯�u���9�{L7[@(2[D�%�T�SbL%���=$�h�N�c�8��6��8����E��&mɯ�E+(�m�,;f},�{��:��LuȄI]���6<�9��B��E�C�{�6����á;�)�C��0����;[�5��a�ȯ�//�Z�)��5S��t��K����GB_C�YS9:��;�mcB�b�tڽz�*��@M����%�8� w����C�cQW*�3�^�.����ap:l��������K�`���ü��҇�o�SWF������8�f�l9Sqs��M���1Q�3(���G��UV��!�	�j0�������{`ܽ�"���#;�pnb����PV��\+T%�N��w�az�Q-Iwz?��m(s���<�O�j�D����}��y�N8TE��	���)˗�G��JJ�3-��	�[�:'G�t.�]��j�楤����}�N��݌��ej�cq�(n8�K����ۥݲ�w�֍��O�����N,�R�F�!6,u�C���f�V���w���v���i[���8����,d�3f�RM>u%��uDPo
��l�6
�|Ta�����:�7,wk7�Q'�T�jg�.�"[al�T�_���d/斘�����7��#��A�e�lu�!�+��Ot^<��C����GJ�����4\���*�hξ��|ŝ����WP���*z�L)�1KXeH!��~|������qu/M���c��ſ,�e���v�+����\ K�'94h����-�Op��dȈ��Y��ۣ? 4.�]��k������6���g-P�9�a�����4vtF��5Ĉ�H�/k�(��*�ΰ����׽��)�G]i}M$�a��Ҽ�"Ĭ
~{���K�ym����CJ�;/�ܨlÍ���x5߳6+C���7h�P�?�6��"�B2����YP��[!�9����'�#x��ͻx
>��(�[I��9Z��R�(��)w�?����-c}�#�~	�Ǘ`�ϵ��P�8P$5<w��>�{���'Z�P�e7of�xE+c�f�9��?���F ��>��>�<-Z�Q�Q���K?*
[_��u�!B�xɩ�Q�
��)�� ���1��O�f��ͺ�휗����gPg�H?;i?OqӁO�^_~�2�r7�O��Y�Ȑ� A�o��ȭ%�r���a����H\�?�;��U��][࿗�	{�����5D��`�u���������$$.���5��� �s��J����i�����噍���i��^�-.{M�LX�a�m�Gy�(��W6`��.N;��aQn.��-�D���{Y2o���D�\��j�a�)�k�w�fO����ػۢ�.v�,�ީ�Yi�������Vu��YFâ�?��5.��S���^��_5��F�g�6[!���u�ܬ�4��v:M�J�}5��4�T]x�~�#s���vl��awH83k ���[��J.�y������x�5+��4�AR�I�v�m���\��SNJ!��0���C�~-j"���F6��ID���5E|(�z�E?J�SN��p�B.34�������o�FwL�R��Z�i��g66Մ7⛺��hH\����=;Z�x��MI� m��<?���i&���gֈ��i[���� �Gk�,-l�V\!����ͪ���;��{0�+���1��t[��<T+��{.��>!�T���u�9� Eh>Ye�7ཀ�ڡ�8@5ir��
vjg4�����S'��S�J ?���$!J6�=z��~�PGe��?���5��ZV�;�k@�"��:=Kׁ��-�^�L���9��*�۽��z���������:����f��HB^�oтO�)m�m�!$J\�]�f�#Z�̨��2��t�Ԧ��Py�۴�ڈ�*���ԕ��J%(@lv8S�&��
j�`PS����Z����a��.�>�0�� L�w�VŻ���o����d�Qd��k �Y���<�K�a-H�΍^	m2�(`oNxQ�^Ӳ���N�"�^g\��IQ���$��/�]�8��4���B�Qn����o1����Pf�E�>�X#��)���n.�>>g>5��G�%j8�5+_�ӟ�L����u������i����6vX5,���鮶V�9$��N�Yi엽_MUm�5��A� �1��Sݣ�n|Ѭ����w�jA�+���#qx�9�C���!]�C������8�8ST�:���BSC�N��[:1Vj�#�`��w��<��k^�c����2�: %(^�l�C�U8�2��	x=v�T�7�g���KlV�K�juN=��g :[�"��nOa	s��7�?-u����Y��g*���ΰ1��I���L���1Qe(�c��w�%h�"e��ʦr|ù��*�A:1����lv�'|��2�	
���l~V�=?+�#�g��"b^sg'���M16�[����a؞�*�Tb�LD�-��(3lm5C	Y�ۛ�_�.���mQ��"���Ӣn�.�>
+��������\̴t'��D�=��G�-�?��������*�:t��+aX���N�N���H����ۮM"D����%�a����C��U��=Yݼ����'�[Y~�F�3}U�^��E�w$jҕն���U?J���i�<>�������1tY-���l` u�4q�7v]�ޏwHs�nV�\� y:
U#R��M��`�W|�wkMg;���K�rn���6ˤ�M����>P����ǧ���Uu`����v�w����|���\W��c�n(���F?�p�^AHB3<��wzV��ޟV��˦�&�\Q��`ҳ:��l�NT&�6��M#R�@��KI{+2��+�qvL��Т�ֶ�fa0MG� ����9U�W������A�'
eq?J�lVH����`�����SOy��pZ˅���cט�B�x�Chk��`pp�hqR '���ǎ��YH�q���v��r�L���T�C��֢���לӉ4%����/��	B[+'�K�dx�/��g���S-s��F��3���_�/>��15�d��t,�O]�h�wG��&	��	)/��E2��R(��Ru%��s�dgԿ�?|$[��g�278����8�z��Qi�_kܤq��,���#wz�	X�J-�p���!P�ӷ�3	q�PDY�_� ��+Na��.�K�m�)�?��u�=�0W��к���s����k@-������YZ٫n�Ӳ�rj�ۑty�B�ma�X�W�XA���}۹B�>�4���F�	u��*�x"|��)�G�wS��.P�]����ԕ�������ym;)>�3�[���$>R�31*џ|;׻���CYĳ��H�H��>#y%�C��=���mP^ �ҫ�K�.n������_5�z
�Z�F[��c��"�Q�_c��)?�F;Wn(���<�./�g�YfIDߒ'��7x=�SO
">^]j�)n�����e۸}�3�%ܙ$�����Hz�1�K���T<P�� ��B�T�d��L/5�d��e���a.���Ċy�o�T��S(���#��Ƅ�O���!�~��A��c�}�"D�z��@�Y ��l`2@�|��I�j�Ә��zͬ�H��
���4�u&2���/(��nW&�YZJ����q�1�m9�~��>����	��5��(%�R�ysRǲ9wvv�`��;��ц��5�,�HD�Lx�n�B	/���!x�þ7�۽�|c0��UxJ3�.i�O5e���:XܾM�fa�<S�ƴ�2�l�������7!��/���%����o���g���p|d�S�u��c�%�gb�Qp/u�~�\��y�M�g�o"�F)��.ۨ��8�3zp�MoV�JRĳ�eѹ�A�*3����`�� 3�~Ŗ����C|����t�Nv�i�tV+ix)ᵵ�2CV��e��օ�né���u]G~��o��u�Yǒ3�fF�8������=���:���������4���_D�K�	�Tl:r��ĺ}RԻ�oC��h����3������p�%�,�L0����E�D�0���-�HX��pN I`6���*�{�y���w����3QUƔ��S�p�`+�O��m��Y�'��p)^|�G��p_**��d0r���P��N�2��ɡ�S``�ela�G�n���#���R��`����@z��;ӛO=7�1��~����r���>!��&����W�f5'İ
	�q��VE_T�{� ��4���S�A�����;ęp��c"������K��Fe�=�+�� �$����^�v�W�`�>������潊���%K�02�Tu�|�p�Qu�|*�c�3�& F���Ža��m`��`��L�I�qS���`m�iy�*�g�оU��| SP�.*��%�ӳ{9{��1�;��s�j��{�V&�Z+���?k�������A���m��	s)	H
��"j�*QIȿ��;��#�[�Y�4��{�ѧ�W$R@x+We��i4$sn��viD&��v��E~�/�y�$2�~~����|�R�A�_���� |�*���eg�՚��n�,��| ��6*m%�MR���
��$�%q����d�Q(_��⠗�׉Z��۩$&���z+x��N�}���+5rU���u�w�_~�����/Th�*n�9���'�Y���i$w�>�����΃�o�J=����E@��4�wi�?�7�)Z�M�eq�� ��	�!���x`�ax�j�EG��u .�oڒ�˪\�yv�F���N� 	�[`~����E�Қ���1��Y@v�d1�����%�/i�k��?�{�T��kK�mv3֙���F�����7J� s��l���;HGj�7�K��������tʈ�sO�D;�窙8Q�����?�e��D�
�͐7�k:Z�0���|��-G��������@f�~3zA)�O�4a�;Ƕ��!�\�UW.��ej�����9�YǊs|�9��;'U�M������1X	�M/L�]߰�[���o��>������4�)��3��~�O��������HB�5M���,`���bF��H��5����;���IW����=��;:#�>��Q��I��<g��[oP��a�֤4c$�q/��ZS�%-Oe�Z�ƿ�8}��g�t}E�a9,@����M���?�H�Getǎ�{�q��@�ُ{��f����m�wM�6����'� uȚ��"Р����i���w3�7%R͒�[��+��O:7��q�'>#��=��:�d_,4y��J�
�6_�R�I²��T�l��pAʗd�S��.+�}=�)6��7�Y�0h����>��1�&<n�B��qw�iK
<z�&`�v�񔳧�#1lȳ�0yZ\�l�;sI)��.�2BS狽X$r��u��B��a|C����/�����y�[�**ym�����E3�L����h�i�|{�|0��F)Ü��r�P� O��;[�M�흲�i.���*N�qA�L��MHN���|���0n�p��k2+�=��RR�p��v���&s�
FyIq�$�i�Oj�PJ>��Ny�����_�v�2��ۚ��3�>��o 	!�;���*mֽU���
Q�Va���E\[sF�˨�����ub%g�.�����i)<�g2;k��A�������R'����*�m�l	���'PR�jND;<�&�f���󴻧���ʷ��)���Y���񌏹z���٠����#K�mȝvg%�j3MAr�+TW]�CE�B\:�N�}ՀLq��پ#O�{d��k�܏
Pvm�\�f���nn�]ôB�.��g�YƤ"�����K^22�KR���e�8��a�_�w�`N]*�x��j�����D���w7�{`��ʼ�yO��������!���z2����F� ��}�E�Zː���t���Ӱ=�i�n.��2`Y]
r,�6��I����ˠ�d�ѪtuH�.�å����X����;r��d�T�7�wV�{�ӑӻw3����7L��O[�a�'�^��\�s���k��Z>y���mɊ��P�8�+ܷP��� ��6��l���`30`d�5��ߓ�� �#������� ќ�1p��D�_���Nj�\|:��Yz��k_�~���1)���6�������'ꤑU�)�3(�aD��q�g�:X�`�_��u,�-l�� ��iM-�<g:�|�WRp���Eˈ)3�v�`��\l�I'9EM��yM��[^Q;�ha��F<h�G.$U�G���.���8_�ž+��Snj��]=�V����>G|=G��N�k�_��nuT�;k�_j]z��dy�V)^u*Tu�۰�����,_7�a��N#��<عf<�r��� ?�=�Я��_�V�bV�:�u�ir����ä���E�u��� ��Z��?��@ΨP3��0h'@xd�d����l�U������������{ ��ߓ;�s;%�꼢5
}MN�?��=����P[ּ�`tG��/!����}%w��$�N����DO�2ËgD�3z@_[�4���y���jw�Lu�x�ܠ��0�[�8G�$�i�|���=r��爰f��h���vs�hD���.�xWo�Z��#��A���j��{��t�W���U�
�W}!krc6Z��3�ji7���&�V'Fķ[:
8;t���(���x*�:p�J:��V%Y���Q�y�yJ�"���R[f)��U����ј\g1v9r�k��TNQC�hH �v@t�l\�� F6��������I��;n%�n|tT���8�aZc|׎G��Vw�9���c�:Sb�u�KPA�<���d_�f�%�*�a5�����j��k<��������b4���_�΂l��أ�$­�u���3W��5G켊��ރ7�u�/��Q5!1 K˶kj��q�s�G�_���]�����3�e�Pg�A�'T��0��W�
R�W@x_��d�W�*J.T�P��{f`4�2e&����'Y� "��������՟�����t�s�C��������0�Hi_��(��{(A��2�V^Mȿ{��Z��!��޷����A�����g6]�CAJp;5�w��������<Eԃi�b��z� �Jr.jec٥��q�KDbקB����n:"��_������LZ'���v�w����z)�bd{�)�5���N�jg���_p�n��A���x�r<��RE�x��$���z��=��yQMk�����w���@NCi㎮��[:�Os��
�������2�`꫄QF�	=����IC�����s'���j�� |2�ɺ؛�$"D%�E}�ll.����¼0�w�<���6XO��(�-rDQ�=h�s�-v�W_�c�T9�jQT�5�l����O�2�B!v}���Xk��Զ��c�q���_9�+%Y�\t�9P�˪�m�lTI��&�qGL���j���6��¦tDP����ڽ�?��<L:�I�Է�j��oBu���@ ע���?��`�7���k�91@�3Q�Q��y���7�ئ�����+��#�D��4��ƺS�x�A/�@��+c�3���K�F�&��-���O|�(�Ձ�Ҡ��V��"�o1�T$o�jM���E����7�T��Q�c��#���w +T�?`�[���y�C�Z�����Sz��^R҉��?l��	�/I1A?7��Qt��i5��U����%`��㻌��V���q�΄/¦�}}V����{��;�C��J$�������(�e��"e����q�V��d����D��J!�HO�N�'Ա,�̺,ٵ�f14op����*�!�pcF���ŃkyO��UQy��ͮ�F��.��BK��Dl<���>j�cd9+gW5m�"��fl�wK��=��m����Y�ʶ"�
L��\S��I_��rh-�/�b�Fm�S��/.��Wld�{˹�i�~�	��V���=ۺ�X?�Æ����:�L�!3�wj�����*�BK�֬�hRs����e(i���W]Ew@\��������v�|��nZqS�985����1���[�K\(Qĩ�����)�֗�W�X��=��7��m�ˏ�Nq��t�i��k��0eƺ3�&��5��Z���Mf	e#(^�3�H�Z'yk������3��|��bDo�EE��6Ç>=������&��*h ��/�V�`1>ۀرk+�נh4jT�> v�)�b����[�[s���Y!����ogk���ߖ��`�}�z�-~y߫�Ϡ�U��)~��֗4�}��_lYZ�vo��k_3��	^��Ăٳ�N�w�r�t�o"}�-o�d}Ŧ$0�9�0�IMx�9a���䙡�Z��!P� y�+d��4rS$��it�h�Z��7 �,w�Bh��º��w�-�'ڕ��1��:�@�������"���[�5�����9��Z���8��8~ߘ`E�"WV�Sy�����_9�c`W���'����7�S� {�*2��N3�\���֬�SNR܅�������Py���G³<����|e���3!�]��C�
�u�@}_~V��ʯ����KVV|�{sGɈ�?ø7��K���0r��n�Uc��!�1q9GU��35�ӡ��%��#/��>�:}��ْ�.�%7��F:B�ʻi �Mn0Fy#�����ɳ:�sM{�0���������c1��]���GBb�ƨ�[�ϻm1䱔[1�����	<�8�~���on+�E�MU3.����zڮ�8n�3�N5�>n�1�N�Ɓ2#H	����������Cp����i�붥�V�]T���m\*�/����;K��k�u�LV�o��ԜMU'�D�݇5����L�iM��xp� o{Y2jqK�D��X�p���&��(�����?���"�X�,K� QvB��B̖�Y���3j˅+�B�'�TP�+�B�Z�O�C"�L�H�>�` :�U���{�TX��o�H�3_}	�|�nE1���Y�JU���_�`~��w��2{
c7V�`v<��ּ�J����l�(9]�o:1�0��\q��v�_Y�������d޻��J=����s��QW�d�j�k��6�V�e�s�F"��z��/'�ɝ����ŕ�&ↂ.�0֏}���ܴz�r���3�8^�����=�����H�=B�/��@n�9ޘ>�!�e�ޏBG��S'x`Uj�=,��AZ��%E�W:.߫4�et�V���3���)��xW�J%�r��M�P��Z YV��Y-��y�S��	�&.��p�?M�Q��P|i�B�T�/tf�k��>�[.7XG�1y�9�����}���i=��#+u���Z:ߕm/�xZ�D=X��4�v6��i�NU�e���` �b��G��T��ӊ��{W�XQ|^�p:���O�ҹ�-�e�~sҪ�鯸����銱)�Wc.�����X�G$��(�ιCqs��I�<Įj^jd���b�x���wC+�'A������(`����um�o��h�iSՑ�cO�PYt��SdM��>�*:��E��O�f1�s��1�7�^���l�dU���,�\.��G��d3p�f�jڌ�x*[`uJ�S�v��]PM]����L?a������F毠�e�JGU��X����Y����z�mB��zKsӐ�ܸ���JN��!���Q	��'4�[w3��[���e��޽��'�[�_Yj���Xf��7�F���R�(p�q��I���z�����
�v7�i]_7Ae��4�!|f	L�����1Q�}��Y�I�#?O� ���q��׫G��)���i87�0��$W�_;#��R�
z��]�\� �}���ZP�4�������nf��XV�w��)����F>kX��s=�,�9�(�o:{�ӗx����}����"���e�ڇ���C�Όu�S�^r���+O� �~�c��0b1�v@���*�I��7�.6�)c,�S��gR���E��/$D҄ޕi��ێ����3L�߼�wz���E���&jT�f��z���k���KH-6J����W#�S��)(o�$[̚7X
oL|,�s5�Y\O��ܳ�
M�\���b�ύ�a߃�#E=��!���=�)2[����^/9���S���\�c��UF��4�B�'������@u������t&g]rH�I?첤/dG�THm��c'�fԧ�FA���Yd'��-�8��J�2�h�$��h� �#c�Ym#�"B���K=���Ry�"��s�+��p��/�p���b鍄�k�,.��׬����q�g �w)�ї��!Tp�9�t�T���%���^[3'�Wg[�?pAˤ�-���V:Y�b�_�9�lZ��3-�u�M�l"�a��ֽ"��LG�+���͌��?��C��#*��Q��'���w(�P�vܑ���%�U�Z���]M�{�e��[���8�9�7n�����yrW��;���A~���oB�0`A�I��a#��3e�;8Ů�|�t�m�}�	P��>��4����
��J���]�V�R��حѬ+8� n�2�lv��%��oY��y_uY�b�'�;*�"k{E���A�G���������m?/9~�`��J}1�͎$Yv�r(̞�Ң�����f�Y������߉�<C7�@�Q�Xi��,�y9�n��S��p۰���,��f��t*CFS�xK{P�l�#f�>1�2|�鬂�|�A%�)ǂM�S��b�� ��ڂ�
�|�ģ�!���茄�3F�����Ґ#+?���F�u�1Rd�Z;�������;i�Sc�S�.�7�M�r�����g)������O�M�l�oƂB�[�'G�2L;�U0k��5��`��L-m��#X/�2����n�q�����s � �Yh��0�֧8��M���%��`@[+ڽ���j)�K)�g"�2�TܛQ'�Q�8�vz�SR�QdMM���Hu��;۪.K3�����{J%���	��9/���.��ԅ�P�����0�J̲�Kؕ)Dx���萑�Ƙ8�E�'�.��{�H�(����k�x�x�g�����;�s��
ͥ�]��t�f[#�:�]"����6"3��b?"�λ��� 2�)��m��+�F~>K�F�3v0o2�]R�����L�B�ЉɁ�����&
����ܭ���i
����]5\�R���9�0�����KfH��Ս@����u�vP�!	NPU����-�\Z��G� ��:�J���q��
�){r�Q����{p��&�N|�%������m���������;CP		5�gM�U|�O)���<2���4�V<ߟ��W��+�F�t��ޛ�+W�1�!��irNܢ<2�_��+����4�����Q�z�6��d�#��(�S��`2[<D���/��>��|5"9'�M�3������,���f�כuG����:�W�z���Cj�����kb�ɰ����w��۹z��{��ٌ�k�՘�D2�^��"���\[����eL�>���rl�	F�f<kD�m�I������ߞ�oZV�'�f�y��s@�T�mW���@ J�_d��q��i&����sh<�f �u�t�cK�S��i������|z	�� �;簃as�����\R�ztì��Y�t[$G0��.y���YUd+If߉��U�^Jѹ�-�����0���l^�JX�@\�Ǝ�烴��ͳB���a��F���Y��4@��].߼�e2�rdja���Q�3���kr�O?ra�W�9!�V��������\0К�ш�p��d�HGP���JRO|fi��\��4d���b�&2��:�F�	>����U�l�lf�Ȧ߮:�Ca'&7L3]��2�\��E��YQ���NW� zr]4����5 K
Rp�N�/��@�v/��q̸�.�����Z�Gc�<W���?��eJ_�/��ܰ^�ǰM����{:x[�����~�N��X�\	
��ݔ�:�!j�ƕ�^Z9|��1l �� &G�*�6Dt�$��p��@Y��-*0�犲�HSg�&���7~������	��/���!��s��PuHu��ϙ�й��B�+���|�!Í��C��T۲l�z~���f Mcz�<} �ݿ�+��>�#�+��q&,�)������R�R�4�9�ݽ�jV"�{'̆����m7�'����){�O�.7�;�-�J�܆��y/�+���L�aE1f%O�[7�d������!9e�O����/�E���W��F�ީFT�`O]��^�S�]�TA�*+��N#hD��]��"�!�e�9�.�l�Fy��n,_��!������əOi�W���M�u[Q\���K��n]ۚͰ�s��S�gEev�#������졚���Y��BW>L���o���9\У�-�>A�Z9�=h�ͪa%�����Lg����F앥�0ٳ�^���9]�5�~�TV�x�4`�!>�se5�0�|-�nσ�����2-gX��%H�dܖ�TەZl�tY�-��D��v���қz œ��`�/
 ��J+(�I��Gx2)5�4�8~��n�!�����5�"����<���}cFWܧ:�1:N~����=cqfo����0� ��z�S1+q�Y�H�ל�{\�i5'��;Af���������I��&�n�V$SRh���)�tV�qtr3�j]�tuN�*vyy�Zf��� ��.;X�Q~��E��5~������yp�J��J������c���2�z&�E$�7G0��[j �g�#��N�vҾ�ϊg�t%V��oZI]I�UK�Y4oL���N���I8\<~1����?�"3%�˦l�)f��?���D����ȄO�/z���KD	�6� kf��8o/�`�0~�$m���V�׷�Hm��Ծ�Z�����׏:�,�/k��������y�v��%.���	j���c��XhE��o��I���+�����M�?,۲g֙�w�e�Y`S[J����?�N��|):Y>�����|S��m"�!��7g�V��m U件�����?���LGP&��STۙ�ڵq�\F�k�>��?��"Zt��ѶE,\�~�*�u�h��'k�!�p6��sݒtX��޴��(9�8M�WB<�5���d��s�Mkr���Sm�/�f���nv��8��Cp6��,�N�����Kk�Bs�W�F�L��"il���1C@b��ŵ��8
� g�����i��� �ٍU��)����bb�H���Xuxn��H��>�w٣lo9r�� Qz��sl��PX$�`�MMӊqu��Z�3)5�К����= �I�H����-F%@+��7�pp����O�n�}�h"���{�<B$���<x�z=�u�1�/��呩���thu�W�8A0;��~�>�e�х^��j�����X�y|7c��e��@�K��F飯������J$��x�}�[o�������E,�AQQ�nP)��&!#�:d�ҝ#6%��5Bb�6r�����}���8��s��y��޻��L�po��#�M��"��#_BR��_u�kϫ�Ϸ7J�(ǽu4�^�y_�.�2|Oe�ǵ��/��E�W�`͇hlW�Ȉ�M��~XJ����1Wb*��qR�}�\��@\���\����Z퍆��nj�ԉڥ+U��Nu�c���Ch����!极�8�bƘ�����8 ��fζɃ�����ʋ���Ƀ�G�ubU+�G�8r�H���QS�����h�{k�k�O�?�?ZX��H%�����|Z��H�k�	�d)dF���SI��2$����!	� +�ke�����V�7|���	>ȍ}BL���%��o�{�6q:C���A����5��<H��c��rȜ`v����琯�̠��9�~y)���?��q4h�ˆ�I�/ӽ�J��z�Ǭ��7�4^6`Yf�n����(�[s��<�k��Ik��!쐶ͣ*u|�N�ڝ)2�r�"�N�����;W��tl?�;�6۩�SⅬK�vNC���=Q0�J�q�K-6�q�`:��W�����~�@��sJ$n��话�9`��4�C`c�J�QC�6գdo8�%���D᯻����[�3�J���Ux���G/�̚�8��In!J�D��s�y:E�?��>�I�_����v��tx�z�S���lu�Y��S@�4��Z�%�B����:�����mt�ʧ"l�X�����N��,39�S��L��� �%���=�@�+W�)&��rD�ڸ�9}ϦR������?R�H��u� �i>x;�)�'MB�zB�E�..�.���;ƚK���[�SG?ɼe�46թ��� y�G�ߖ�˳N�ћ���<�~ƉC\4k�1�Q%���! ���^��$����ɆL0�
*M"#�8����gG�-�:d�j�����������Ⱥ�����M_7���냷:R����5w>7J��%3	[�.fL�?Ѳ�I?�YJӈ�
ήb���S��[�5l���2�}<f0� �ͯ����B�Yr���p�]�S�74�٫BB�E�Yū�M]=a8#`�ekv�|�&�'d��9�P�1�BN�n����@�V�ѩΓ����V�i$Ef���;7�w�_��W������ T	b
�1�ݚ�|��	�J��eUi��Bi����B��N�|�(���->���ŕ_�+��c�w��fE�+�S,�'xLڮ\�����r�/S��n�|t��im'���;d��R?K9��N��W�-	ׁS�6�P�n�y/�ʗ��Zc�Y�=1 �Dt�Ovs"U�̃����6�궗��	�,�\&�r�o퇯 �uF�9��H��pM��)8�j3�ԇ��]��z�Ss;��X4J�HM�sQ�S�bcC� FՉ��-�R��ᨄ%��!�T�S�?�>�Qmb���F�5+�Ӟ�T��<
�c��B��\�jH�|4�k���o��館?;�ψ��0["7O�y"7��/�@3�7Ȧ�rb8U/�.�{y�z϶lENI�R��g��~Q���v(B���Y�m��m���,�D
r\∯����'�z.����;}�5�lQ��L�����s����!j����\�9�t�\	3�ie����������j����5�5Ե��F���Yc���d��*�t;Ƣ�Y]�?���*n:�����p����%�)��'!F���U��p�/3%F�o������.��c�N`gZX�nR�lfvnU$pYD0/�V\??�;���S��p+ؾpaJ�j9@�>jes���6�A�d��Юu�iHG����OD�T#��[bCg4F�&͘�U�G�2�5�L��-�"��*��m���Ut�틫�����Ix�se�SD�*�N1�8�i�:��R�]�Q�3� 1\Nb�bc+{�WX1�"g_�~&]?<ܚΔT��B!FS��*.�y<t�.�~ޟФSj���Cs���p�祝�QApNJf1 ��Xm!%#Ο&R������8M��kdDF�qT|��f���ŋ�����\�@@������h��*Y�9�G�8ŷ&�y� �+'n����L�J/�X~y{5�Q����"wD�u���tJ��I�pg� pD*�!�G�{d��d��Lв���"rI�����wg�K-� ��o���f$� 9NDo4�p���%������H�G���_�/"Rv�-HY��v�÷P�aX�Uv$��&�@�>��79�_5��B#3����Ő�/}�FQ���"�e��><�T�e�v�|�r��L�J�C��(ֿ���(��~�����,j���Ҫd? 7�w�0�:l�R��WrO�̢jw2�;�U��\���G2�z�&C_Ԗ;�d�d�q�a���w�a{P*�~�t��:=�	~ �o���zTN��~��w9�@v���Y&Tυ�ߚ����Z����~"Z)��\�	B�6����r{T���O�Җ~)9p"��@@z�$��U��@oURH���~��N������^?��y�F��Χ�'��=���*{���/k@�s�h�{3u�E.R\�����}Y��n����0A2"�p�f�w��R��[Y�*��r�s*�^Q������hO�K��J!x�r�@pc?S!f�^-�4dD�+�GDD���K��(~�:p�W_�#H�s�0ǡs�i�g�؁��o[��+�u��C�h��:���\&�[����kY�ҿ�18*����[bp+�+����vq�|�:���8b�)����M	�DQ���A˒�s��J�j���˄�w�����;#�Uդ�ճ�G�}�aY��C��H8��9���и�_M9~is5p��@OAE(�+����rMZ�CZ�����g��?ǯ�|���rCM��^WPA`���7�`�!��{.��,I����L�L�L^J~�L\_Q�MnMʙ�������ĺ��Wz�򉇔�#ǝ��,c���o�Cv�s_������k{�MK��P�>�����h�h�	G�:�+9�~5l�#_���}�~H+n��7i`V�mm�ep#گ�L�(	H��J���ɟ[pt-u���� �!qY�z���lU��]܋w6u}��e�>>��������l�$��ex���?�o)WO�S�<��HF��t�۱�$�旡��m�R��׍F�Z���~�x�7�?�@&%��r4���V��iur\���PF��u�x�P�����{�F'������JI�3�G`:�w�f3=�@�E��%M�j��UՌ��������9� 3����haTNڏF��9�<�RS�3������%^w���/���Ì��x���X}��ʬBS�*,�(,����̔�$�
�7���ϴ�n�V3��|�G�\)ܓ%l�h���O��D�9�?���Q��8J���-@<���7`�7�b`��`ݰ���F?4-Tn�g����(}4����� ����7�ʂ9�{\��<������	y���m\�ۥ1�F\��W������z�2+\MPe�����--�f�U�X����J�W��,���U���w~.B����~_���V�;o̾��d����xC��3/����r���4�h�k-O5��&��5���h�I7��J���n�����!��mkv["���^��|j�"�GC �w��Y�u���I����T��C9��l;�k��{K�<�[>���|��R3~�Z��=�j)�c���_���G����2Q������?���MF&���'iH�m҇k��݄�c.϶���-��/�k�-���v�\y&�y�� ��~�1ۚ��
ƟB����>��� �!o#DH�-=��>|�V��#��8��i���G��o8�O)��J�v��{��R�[�%�y�:/gWX� {.��p,���Y��z�4u�ca"���]C�Vwed���Le�#U�Y�G.u1o��|���1���ˠD�� J�*�?�eM�_��	�o�U=��,A�:�c�O���l)�����<E��HW����\�O`.,r�Y����ϵ �C'35a%��/��I$���/����꟮����n	���u�Nc�,���"ot|#6��&�7�W��W�s�âT����DH�}$vM^&X���P���)h��IO�o�l���4�ܰ�&BP\��uw�u(؁��LknBZ���Hqd����Jx#|�8�;�KIB�HX�wܜh�{!�,�	���ԣ�v�x����U&�(���t<H.C|^�	�������^S��tޟ������F-b�'��m��N����Ph$�K'�̿0��1�/HS3]�t$U�/�]��|
��7�e��ل�®�T��,��U�ڳ0�G�N�92��'�M�' 0��Lk�T�4�]��j���&�߼�W���B��o�k���.��!��Z�#���Р���/�Hp��m�����'/�}E~����t�ooBʈ����3�&���X�Uv~�8�h��T�t��e%���؀�����A��	�٪]�y95��g&W��U�j���0��@��şjTe��cìG���o�7)Q-�ؗL2?��}�=�PxF�&2ٲ�q
u9��m2�^��+2����k�ը�����^�P�������^�otޱ�� ��|:�]�4f�$ nrg�3F�)�*
�b^Ec��s�Yf+�
�Lε�����T�8w���+�P=���	����K6`U��׉Y�-��7k��=�����~nq�z1�K�����4�N�c��o�3�JC2_��ϔ����"FF�ƶ-E%����ְ:�����Δ��= c�1۲�8vJ⛥ii0>v���&�7��7����;�e���O��v�a�r+�B��\��Si�������R�������:YB9 @F�B� ���%y3���C��Nx<�x�Op�~ �9��{o2��R�kf�V��B�۵� ��,�8E`v4r���f����qX��)���Q�%Wa�����ŚF�pRR�X4@�t�ԅ�7�Dn9-�E8�n*g���v���Vw-������V�̢�̋;��4��"x���aY�6��L>���t���[En>�oPv{v��Qnv̠�q���,�\vC��^d��ZtJ&ǝ�w��]xgC���ٷ��?6*�vs����j��6���q������:�5��F��D�Y�0��ʭ�`B7횄���-�G���d����]����p���,a��8�����/4�!��2��Z�����!w�$�O�����M�)�4]��{� ����ɔʉM������'z\@�t��M��=�],���h��Gr�s%ݜLvu<"Z�(^c�3[��i^f��px���U惀�O��+`8ʗul,�y7�6� "�C�r����cN#�b(ZJ���$����[�l���;7��v!��/��y�n��ն�K.1_���Qʃy�Rw�����R�J�\�����O:��iI��[(@Ë���0��ĂNk=M��Ѵ�Y<���Ľ��9m��b>��L�{���U�!��)����$�������T�J(�u`y��Xm�(���v�6f}N���4?@�Z�=j��B?��ضB�����A��X��v��+���}?��H�"�P�#sI�/rS���F9Ъ�}#��LhM�hs�)>���f^~�(�T#[��#�}C�=��~&|_�:>Zjkp����H�/|l�}�U:K�bd��9Qu?�0��5r�;�P�H��"�USR���}���
���<�LE!�79�#��15��`\dq3�����"T�%��4�����I���<���J�Y�^}��#����0�%Y���Pf��@�2��GtA&f��M69-�}���}h��P�+e5���6�e�Y�#�lj�J�RS�e�d(�Vd��ϢH�d�8[6zp��w4&���1�_��?n��_?�4�9"ZA���B�������p��F��-��UR��(�̦�0��ڪ��y�F9�+w���= ���yy��I:�֬4��dqR���!gwu����6ã� x����l��2x}8��ܷJ��m��[����"W5��F<r�#��0i��FN�l��+G��7V�m��va�)¯�T�N;�fz�-�_�VK���ʵ��V�r+�F1�GC �b�	�4���D���Pt.aC���b�Ǡ� 9d��È�n�_��Z�������6�=*9;��	��o�2Ί ��i�9Id]S�6��\T?���ea��Zh�e�m��9�W-��t�L���o4����B]f�B���eQ�[�M2"�'�R�Rqgל���%�����j%򵴎�6Wov� Nx��q�"�f�:�v�ʭ:�u�Xi�K����a�C5�):��T��O������]-)F�"9I�'���2�b�;ƄL����ߡ�^��I��V;��5�BEf��%;.����TNT�n{Q;V ������@�e�#M����N��(;b���eU��7�49wr��#XAs����nٓ󺎗���R����pKAR�Y�i��[�K�K�! �����Čs	A��������p��r�\pS�~�����j�����N��X��ȪN�����ڳ)�_�
A�c� VE��fY=��iE�O�59�C^�0?��'�S�r�6o�d�?�G:�H�)5i�W�����[^&�89����x]�/[0�<�S̒�߸-+OU��\^wh����Z�{�}8y�����y�K�]���m��:�J�URB"Ap�^]l7�3ߗ/��l��P���3'\�������7��\۬�v�~���2��g��`c9̷�]i�J�>k�&�Se���+�*=��KN�8��hZ3.�6��&�n�]��b��J���z�c��/��N����?F��C�ٺ���1�|y�_ܜ�|64}
����r���>(�E���	+��o�V�v�Dqo���28����?��{�у�\�׹TM�Γ��}z��>V�i�aX~�$��w����Ss�^��L�߭u����!-���߆iDvj�W�M�W�ǁ2�S����Ž_�I���
®�5�O~z��_9X� �O�n4�կ� X�\� �EnoU��K���3���m ɴ���xǁ��=��:�ʶ�2 '���S��!y��,��N�a�maU�1JO5�f�Pؙ�p�\�-�ֆ��mH���kͱ�>C����yռz��V�z{�sd�{��49�iL��? �Ku �i�|��9���r����|���@$W4)<�ݴ;f6�:�����|��e�=;�ȥ���[��E#.��lo�{H��WO!�[eJ���-�e:2"ͬu<5��Ǜ���Y�\��>i?~?���po�n���Ї��C>�%�_���h��{�󝍮�Kb���/� JAs����G@��0!�k���Jnf۸����{o���ع!l��V�{���}4���H����*N����΀L)0���c�7/�<��2��(eR���UWb��O�h��{3�a��[+�l����6�N�5cShX�d2؎���ZQM58���]�}�D~���%����S��ɛ­�pe;�W��9��6�������_ɒ�0I�K���V�h\T:j �E6o�i 9=I|�.0h.ۺ�^c��`tf#�bBI�x=��������a�P�y��lM�s<����E���{&r\��=��*��9�N����N�y�o��ZVd[3�[[m�:��p����N/(�c�Z��p	�d�|U��:�:"�I~�J��Ǩ��3����/=F��JV^�>M�����IPq^���6�5C0q����&t����T�_�����5�1�O`���kwz_�2Ɖ�_�F��Jn���L�����M�L�s��݊�#XcAo��h�j��/0�(A|�_�j^�:{Lʚd�z�r�,�(}��bo~���ね�Ge�o��r�{4����k-�jqs4���T8j�g�;�=im[��t��}��d���v�p����zu����8ҰMҢ���Hz�߷�%眳��Q���/�<n/��Ҁ9	�M_��}˯>C����M��t���W��<�^���Pu&(��7��p#;�{�唦^R~/g-�l��^� ȯ�N��927g=���F�N�ӳ��R���[@o��ª���K��B��:*;��u��<2��1VG�(��Ŭ_�5,C��T���~6Ee2�����p8����ٺT��^.������K;`$j9!h�ѐ%������\@���P�,"��VW���۸�B�th�}��H' �K�;����N��:o�'��?w<X}�t_�a��]����u_�P����*bL�E��2�Z\�N?Z�8����/Ff+����
$�O�"����Z�IE��zi�P�z�z�6��O0��'��/H�k[<�x��Ŗ)�1	G`���^��qd&0��72I(���X���h 0�6	'�|����F�oB8~VDJ[�#�p��6z�3�h���O��O J1��'h�*��@f�x�u;��@�I�|[�C\?�/Cձ"Ԥ�Hͫ/7����k��"FK�n��W�J�C=
�3gTTj,fNM*������8Ko����gW^<g�Nݹaxj�"-�j���
O�x�5^��|o
'h�G��^4ى��L%t�_���%"��hSȑ�ϔ��������T`���.U���0�"I~�Hܵd�z����1l&��j���W�[��{��-I5.b�l.����j�֯>V~"���3�8�ȏ�✥}լ.�3aP-ˈS�|��y���T�Lo2���t��@ܼp�a��2+�1�L���З������0}>��(�M�3ɩJ�����A��78~�A._0*�t9�#*`�S����N�/V���#��d-W`7,^��2���}�c~>C���T�}{���>7`���� ����=�s��BI*QNa��l3/��jN���@Ff7�ٷ銭�w���_F3��D!IE�E�.��>a�g��) �e�2���[���R�wӽ��>�fY���<g��z���߼V�Ni!*l�6�t,AƪeͲSc�C��~��f���պ�����6*<�6�'ɨZ�r���Ő�]@�Y֎	g�Q숰{ �V*,V�3x���`#Z���wyN��m��>P�[@#��Zŭ�[��R�f�+L�;�Ti�:2|��� M��/�|�!U�g�M��_�-�\����I������i�?1u�ʢ>͍l �r⨾־��%�S�^[���_4G����Zz�y�;��ka���3}����Ȭbh$hQ�Yq��L��ei B�sK9������E�=�V{��o>-�
� ���F�l_v�o���ž�m�A�c�k�\�%�.c.�m�X"�� �>��A%��H�	�;sb7�^`y�I�jyZg��2���(xΝ����Y�p\H@9��=٧L�xϗٞ�3�_V̩��ه���%���|z\1Y��s�<��x��g��_��}�}���t� ������ߔl�671��P�� �����v��xO���D�5��r�;Ǆ~!rc�8߻=!��U���H8��̝����ͱ�Ά���te�7�F,�,������}���o�V�]��s�-��;pc�n)ŬH��*�����xX@�wn߸��*��=`���%��C)b���32�x��}�����y�{���<\�2-Y@�R�`����i�V��5ĉ��=��ޓ�Ϥ�SF��l{\��G����o0�*�����Vƚ��&f�R��t��P��1��D��������;�(�+�+n�)aYf$����wn�l�tރz*��(��	����_]a�a��H�9��-{l�Ȕ�'�:�>T~� a٪H�.������&w���12%x���m�����ÔA�,ȨZ���&b��_Dr�=���MD�� ޫ�+ºp�����0�m��ul*��ꚹhhPP�Il��EN>���a�Vg>��쪌�?��������I��5�A}��f�Pv��m�i�uwܡB_��I�C9�5`�*ﯡ)�m���ŀ��Ï�������x�N���KL������%\z��qF#���N=S�6��z����s��r��d,�H,m8s���I|z���$��|���޹]��q�+A�����5�i�:x:2"F����P�l5�I�ǵ@^���З\0ۜ�p�,}J٩�qM�K�
P`ԃ߲4%]�Ox���繉��%N����ҏtm��<��+��[ps{�ȷ,� I�Gx��3(%�%`��
=�c��4# �!�e�������6_c!�=�y�Se�$r�k�'oO"���
�+Q&D�^Q����xM�7�Ĵc����ODc�a���D�������b�H���;�8�!���@�H�6�]?do��g� ʌ_���pih�$`����:!=���A~�o�	)��QET�7�v���<��E��U ��V��_���{؍M��5-̅c�ܑ:�� qώɠ87`棙�WD؅�Ua�U���R8F%��w՛��q%\����++j��]��
l�R��N��ӗ<�W���]TsK� ���?ʎ��=�X�l�&U�]/�MjH�'�
�"&F9@�p�����8°)�h�P��J~Q�L^�7����6o�/�r\-a��(0D���� l���۞���ݕ�wk�H6�!��3�=����D�V���c��p���ᕈ��G�L�����ŃrmJ:�>��/��N��X{9W�.4]O���2S��t��6<��t��qNF͞[Q#��-���ޕsD��D��U�Z�d4W��_s�W]�N�|��)� |�8���u[Y=
���S(&���Ig\��F9�:��G�SՂ�Q�(�K���5=��k����z_�E_�����&�#��C��XT1[��/c�*n�������7J{I��n�ulP�,��F,��OJ��݆;��[��x/y���E�J�_)�{���+ �al�=ʱ�O��(i�_�����S�bi�q�Y��[������g�We�Wn�������`��.
����`�P�M�h�o�,�'��w�Wl��NS�� �]�|dp?]�����H���;�k�$���i��D9�yĚ������/����c��5Ҧ���F�C$�k�zѧ��#�5Sݪa;-��TK�WW�BmNt��e`�?����}����#e��5�p/Xsh���O��V�[���s���Pcp�7��8��A���J��R�9�#���0�ۣ��s=��b�,��UTZ����@6|"_ ��'6$�mv�8��e�i�w5K��*B�f;�]��Y���@��[{�d�	B�V�%ڠ�U����m���^o-TNl���	@����p�V!̘W��5�i��d�?��A���}F)?2�bJ�:��[�2!\X�Nr��劉�n�`VO�*��/�U=Q,�C�J-č4����0|�OH�v{M��jh򆇎3�]�����ӻŇ��x0�pW!q�u|[w�a=X���+vS[9�Wž�xcjF���	�������а�Z�y�nEe�Mۙ���฾�O	q�ps��x�I�i�#�v^����M��U�E|��j�x�Q�����1���MI^K;;����z���4�Cr��މ��:��<qx��|�^(�Z�,;h�jĀ:u2���s8M��"s&L$r?KZ��:�Zak�ZQ�<~���s#S����'�"d��ޅ\î�;�!�롂��0Rf�x�Bf��_�c��D�vMFM����ťQ_����m*�7@9G��=��[
++:�v$�~�)�D�~�zim-�����M�Կ�yH�d���6���2S���uC"��5���*vξ=��G�N���&��T�\~��mI%���''gǭ�o�:ȳ"�ȷa�~���Ο-,�ޚ��pJG7��3���|Eo��6��g�<���2�M\^}�mx���<���<��ہ#0"W��v���{�Բ�V?��X#z?����Q<�*�C�^�}��͆(U:�k"�;Q��8g�>���Bo5<ΖL|3)j�r8���k���L�Sp��u���4�U?���. ���$�p�'��\��M_o�[G�ס~�F�!�8�o����{AX��b�|0�)�+PLq̘�ۄ� ��W�JC���P�.Nw��cÕ�[)R������#j3;��|�jHǪ��#}��_����_���p��� g���|�n_��q����X#1�U������;���u3$		��&u��.x�G���uQ���Q�M�j����D[X�����K�l��(�;�F�&)ɫCU�i���˫�6��j)Ш7��$Ie-fQ�<&��;�6n��佪�zM�Z��?4h�fB�{��z%f�Y���~�F[$���R^g�<>����|���-?�t�2�J���mJ����h�K&��J�|�0��b��7�y��k�`}1�f��N�6\��!,Ck��ŭ�H�t�T��<���=m���:;�>Q�D~9�]�0&+���3������;�ڷ��փ޲�İc�G�)�WA�����+c3��p��2�GnoJu/�>�s
x�ђ��iwἰRV��D���p�p���D�/�\��:�&y}�y�c �1�c��%s�uثХj� �E�E\2k��]qܓ;�TU��/������;��i��E�6�/�-y��ɵn�B��wy��?��� ,�He�ٝw\�ϩ���z�g9X�&���\��uKUYb�ǯ|v��1�57�o�;2r���M��t��ޑ���K�nN,n���~Jva�ټ'~��C���(J�H`�L�}�tL�:��!�k|I�Oj�j-a���`Õ9����4^��3|3&��j���0='�ѥ-�y��(��ZH
���4��?=�g�ũ�/�.a���5.�@,I�"q��((#^W݃��y�/�4�@|0��(t�m����{f��e�%6``؀k��u�R3�N5`x��\|d�8�]�C"�K�u��؉T���ݎ��{aϘ6`r��W��$�F�Ϋ����'i0K=��A8e�^J�H""V��1��2�/R H�Q�YWO<>Z�d7`��_�
�yƃʗ�DV~
-W+9r�C�0=��[����tf�>j���q:A�]r��{���������3�����Ȓ0���j<~�v=O�z�3{��x�����{�`I���M�Zu�+"7_�����>9��~�`s�d���_�������죝�D�qII�]
�?Q�n��,��KG����.[����?�i��oT�:�+��-w؟��"�ȡ�{?�]������v}��zDҡ������~t�'g�P�k{m���#'M���k���4$
��å�>)���q2`g�/	��o!�.���Ve��0���Ua�`�	�Q�IC��s��)�UĐx��"y�Q�(O3!h���ȿ%Oh×�?�����T8�����'�-�$������9��V'Hr��������[�ј�j���� jj�#V������<)ZP��m3��9���8����qi�)��1�����s���w�X�͆�[α|���N��>0�+����m^���cՐ�"rg�;��6�'�~�P<�����O�.Ь�Cӹ�"��^f�>J6����;�É!'o��~OdaU�@n�����(GXq��Me��&x|9��Xw��N�~���?�G.�,�z�et����*��sP��tk�W�xǠ���s��ږ�8�ZE�&�s-�3�up�Y�?��63�p�ٞA{K_�_�@�w�lNMi���=y|�]��=q���W���{�E|/������j\�+�͏�l��׍j�&;�/�)�ڪ��'��,z>H,V����Ik�����-��OWp=�36%T"�[V�h*�l��8�D�R{��ÜM�@mTc|�c�D��{8�w���t3G�
�f�A}��?�<\���$��������]��i�P�c�$��_��O����j8٪1�^|o���)� U���^��7.R��>4������f�X�������T�-��Z�'�&1��;���ɘSN�x�W]���>��;��z�a�_6.8���>�:���a����d��OW�6=��3��
e�D�K]��������98 m@hb �x��Ѻ�u3l�ְk�/# % ��U������Ӓj�Ǽ�4"w��@�N�����XuU��a���F�:�#�au#���Ou��K<Y�?���5�|H5ݰo��N}wK�U��L����B�t��Ɂ����j�����p�P��A���P)���'eB�[����O>5���QI��>���5�o��x_+C�pB[y��/��Oϰ�52�,�7E㼞��%�����^��;iݕ�(�+�H�w�T���K6m����UTlyM'�p	�+$3ݘQ�}���\���ږn.��y�ʈ���g�w�f�N: 9p%�f�3�,>�~���y�1�Ș��D4�'�ߴ����_��-�`�8���p����:�H��gI	��GO��H%
 Qw������n|�ӹ׊���L��Wr'���<�J"�d/`1�+a{�]/���B�)b���>#�k#�*Š36O���8T�n����e�����έ�(�W�S��5�mR��7t��x�� ���J�v��m҃�u�8U���wIGG�!��g�_Rx"�Oc�\X!�BE�f������F'��˩ec�@���a�ZL`����,���;��c�R9Y6j�ʾ޷����mR�������2�����RGL~�:������)ͤ��\5E��p!fR�I%�sNAv���Á�c�|#>��y��K%@T�!�\��>p?�\3���f���[,��������=�r�dn7�R��R(�O��EOl|X��ez|��Фwt��Q��ɽ@��8_l�u?�Bp�?+g����"7G  ���޹+4B�9��N�J0�j��W<�t"5�Zճ?F)ޏ�z��{���~����A)����J������b��\̈́	�4>�Ne�����	��|p�k��{'8ݵJ;^���j�:~�ȃ�23پ� �>����Z���-~>=Y܆����H;�����V[Y磌�iu����IIo>���=~E��(M���"���[�j$TkD�:lݠ��2��5s��X����苯(dz�OSYl��S�xV&��n�������;Ɣ5qh���<�nXײ��e}�pƉ�埔�c,Xv���ԗ~�%���)A)��U]�;)�5��σ�9e�[�T;�V��,
�A�nqi��CW^� �`vy���U���kw=�e=�m��G�lִ�B��n]�[G������{�aV�FM'���r�WWQ(���_m�����lPk����!���+����,����<��Uc�L`�1�����[��u�q"���_�ƈ��>�!鋆�+S}�=�"n��H��F��1�[��t�?p�Aٞ��Q���s��9�v�aR�6`.NY��Z�S^��U�8���hLby����d��bjQ�O>���45H��]O1(�mаZ!E�:t�18\��ؚ/��Qے�P�KEF�e{��}y�?�ȹ�su:7�>~�7�%���K�W��L��Ν��9>�8{gYe��ǔ�ؼ���W�۪!4�^�Eu�1�P�a�T�2�N7'���D{�S�J%߱�����P��6����\�(�+ݍ�S��7,�-�L�{�@Y��i��nk,��b�j&V�����[�V�{���|���[�����5w���=�
�` �h�(M����Q;Fu9�$!�҇�f)/�T�@�o��doǲ�8� XO4߇`H,l�a#}ױq�"e[�4�^"��b��]��a��M����)�T��iT�dK��?�;���8��};|HD=Y
HM�1=�7���f�b#%���i
�";�)+"�p�%� �gt�|2���Pdh^��ԁ��q�x�����,o�cm��S�XPc��F�}�~��/S�wҘ2��:�#�Mz���`�(�������,�q�������|����%Z�9��)��vq�K�����\/O����O}�_���M	$*���[����������?<���6�bŘ�A�eo�1"�+��Ēj��#��[�GQE�ͺ=�-@��o����~���;�LO�J�V����)wL�r�K`0�,rR�7s�ȳ;y�@G#!�l&��?�_B�1	-����-�q;�,��P��)�ii)E�-ڱT �p�O��o�U�Y�G��j�!��ڥ�;���Mzz�-��)�����*����|F�@g�����������RqR��ޤ����*���1�pE����9�� h��!x�G���K�p���}�|8�ۋ#䐦��G{����Y&�a<C�U�|�ð��b@��'�<�8�鲈e�v�VI��)��?�}�ks��m��bU���z�=Wm�Cj��u�5"�}�'�y�%��*	�'��p"O���}S�u?��Dƞ��d�3�H)%��B�Y)-�~�߻�/����W������_d���o\wptX�7�r���q73܂�h�};2�$eK|	��UuY��.�y���:������,�iqWxg�I��+V�����m�#1�x'���7�#�(�
j"q��V��нx÷�P��
��i���ix	�70:���'2�{�2h�&1�c�[�0�E`N&�6ְ�?j�앉��hxǈw�J$£���c'�m�>0iTgQ��%�Z�z7��T=:I?�����{uO�X�0za9��:�凿%��p�Ja>�#�I����8��n�6"n�����	vl���K5�*5ty/�-yrA�ܪ�Tc�[�#ñ�5��q��q��N��3��P �Y�F��+�z�Κg����3ˣ����K+&����S�s��ḣ��2�V%�IV|e� �l�s�ܻ�06y,�[��U0����Ыe��yE���Q�nJ�!��30x��u��.�����ީ��_�Z|���P�QQ��� � �R"�-�4J(J!�0tI*%%H���0�ЍHI�C��}~�^_���s���=j�5(��.������(\c5^SF&&w�*��"�/#�6�o����(��f�^�Չ�00v�lОE�}��a����������S���L��5zX��Г�^=�F�|l��+�#j�����$!b:2gџ;��P+�1�4{�%�mkrk�WF�iT�N�*��Nb�ٶs]�s�����cBX��_�}�xv��9�W8��Z\|��Ml8h��qϭ��{�l�팪2w�#�&�|񿞺�z؅�2�:|�?= >�D	uĠ:�8|t���7Ζ��Z2�ٶ���W�3 �۴V,HN�bw�����Z�P���	u;:�l�я/�7��!�h�a'u�'^#m��Gr����=Wj�.��s$3���L���eb����\���Se�h��Y�cO�1tl&�Yqr��^he���s!b�A /�N�)��e�5�>mk��$a�P}�ֲ��/drO�"T:�"����<c]4�?K99#ј�z�)c��hi,�ơ��-JN���R����q����(�1�8}�;Ъ3�O��\	Z#��1d�	e�s�ݪL��mݬ�m��^�	�#�,��1���+ ��!�5\n>곑��S�34i�.}�%�����콱w'8%W$łe�v�&t���7�3\��5�}aL�Ò�@I�!?�Yt(N�p޺,Wq�?���a�{Il�Q�]L�����>-���f�T�/;��u$3�)����~�k�=��pV�7Z9	�d�u���s�#[>!���P[�m=�r��F����T�S��ӶMW_ϙ��I��a|q��o�'�̹ٵ�I��4Q�;cJ��7k��u�B$�M*yV���U��U#�P�ϧ���L��.��pIi��C:��[~��9 ڇ��[���,��V�s����}��l��r�v����;�F�L�Ui���9L�Ϲ5#� ��8���~�����y�Sѿ$V߅��	�l�Mg��{`/š�A�rX�㮳��tx_�Z���R��'�~��l�S���TCk�_�)v����sĬ���E1��M��u��}������A�� ?����[Φ��Vͣ�oF��^����{�,5/;���x´f����O����o�X��*�O��g"QL�������gK����1<�ױ����s��I#�r���NOڈ�4��*�;1���@������l�%�{cm�4�<�<�}F�~}�� t�qQ�B���&&u5
1Û�X���ف���Q��PW��B��T�����#>��(�P["^:���1+�G�4�F�������&P�zQ/�p�=����M��;3���Vûi��:/�;���v����A�h��VKC�%�9J�C�V�����+sg��c;�/��#��{�A�Śih�]��-��o\C�����KN��'��F���?�����2�ly9\�������w�'���3�$o�f;@˭Em\>�]V=�﹵����A�;�b㓸m��ڲ�\d׆�S(��l^�yfo��7n	�8� ���
`ڗ��R����[Ӏ��*��ο	y(�ld�������N�Փ�/����{�>�8��^|8}$=�v�'�"�Mj�@��b,�EL�nI�Pi����x��On*fM~���(���Z����K�qv7��~ǹ;��gn|krU,�<�/�[�5o��;�O��}M"�Q���nw�a">���l��t�x�>�bC��G��Z�U�\��s�����k�����͜?��~�!��i��g>��K�r���:F&^�[B�2�7��54
�	�i����J	8�݆���d���*i'j$ĵeZO�Zj~	�{z6���a�	n�w���u��$��l����iJm���j�
��J�!ވ��i�I.�W�xw��`�{h��?4��v���YFz�M�W�F#�<�&�[�;,S�h�q���]�,s}��4����ߩ~M������'��7l~I{�3�
7ȭ�|�y'�7>a�n�fw���z�L8utB;c��C�$y��5����_����Ts�ZzcY�4{��L{�֘x�&Y�y&h�y���SO���GxV��MXp�B_޻^���C��r}.A&�#��|��Ŝ����rň#T����1��vP�By��$�O揠_�)��������M�_�?����1Y�Y��k����?r^����wOk�^���L�l񷩕r��9v_���`�&��a��`�e�x1#�Pt��ʽa�����8��.�x�����)�G�֣Tԡ-�� $듕Au|�� $^~��ȓ$����?������|/�Zb��(�-��"��9�&�	��'�c�_�h�	�f?�$)j@�pWV(B��F���
�Ю���x��n+GTRx6�5Ο2���3��~����}8T��2�u� "��}�}*A�A��,�}����g6#?��ha�{A�6�a��`5D��Zcy�?�M�f8}��4�ƴ�!a�EУ�2�,��s}�
Z#�`_��s`���w� �N��נs�vAZ~78_WE
�ˇ���_LF���A��cd_"��d���i���ﯳs��A�ɬˤ��=��#m�-vi�掎ͬ��a�ۭ��;����ļ_Cz���������V��7<���E��>����x_�ul�S���LR�K�ɶ!ݼ��㦲������̄��SÖ6>��9���T���[�gd��x�8�&�{��1<۹.y���RB6��c��$���y�p{�c�� B���S����a��UZ"�UdhەK{(yO��%�T/�^�b��v��{4����՞����+�t}^��
��K��oqlS7+7��"+b#*G.Xb�N����ݗ0�:(ט�P����{���6o���>lY�j�5iP��[�	���7��jܛu9kk�P#����z2"�l���������P���Q	yt:�����z-���	{T�-R���?�}��������'�YW���In,�`�z�����l~����������a6m/�����K�."�~�0.코d*�7�{�!ҷ8sL3���BD�&q42WR����
s��{�Y�~��ȲD),O���on��=vXeb���kI��|��e���D��ew�+���#�87"iz��l��\��K��SM��Dl��y�xySMT�uE�4�.�Ӭ�{Գi�ګ��Ɨ�Y��z^���j���y��� ���bs�0�"'-�S��3��ƨ�,��z���s������(�������Wҹ���5){O{����e��-�<���b�,��#���:�����.`y�����!�Ћ3U��z���(�Ь1ص�h%#`��d֍:�x�T�Q�T�����X�����[�I��B��.�f"͂g�FnL�D�m^D��wQ����+�d��-�hک�� �NK|�I~��p��:}W�$�nL �lY�.�i�lBL�<��a������Y��H�P����׾H��7I�塥��>홰��,z�W�hv�-����q-���8��g�9G��<�Jnu��s�t0�>S�"���f�R����3��8^���g��^���`e��p�#�L�Z�p�	��h��O�EW���^K9�R%�YUb�"�j���i�k})���x�2�>6Λ}y�� f]�y���	j��H��\��[�ְ��3�O��IδDc_��D��⾠�q����α ���\�����?"�a|B�Cl���Nv#�磣���k
��ѽq`����ƃ ���H��2ׇwpg(���_;������~K�nوt[}|+U	~r�b��SgfW[%��k�,�X0��gS�)����s�p�m�7�ĎBB"�z̭&��o,�x��pr��8���V��b�:R�N7>~5QjPv�p�j4d'�����F��&�뵦R��jBa4w�O����_R|�t��@P	M�0��>}]�E�up���м+k�3F�x@�>�:��w�*c��kQ��^�HX���rf�_D.D����c�t�%�c_I��!	:�Kd��R0̹+���\n�D�H�3�/�y9��%�軍�nw���l<�=��K����9R��G�s'o�M�zv��܅P��>�� ��a��_;9��[�5�����P����͞��Z
�M5`3��C ␻�͡�-5lK�ȋ�����ʼV���ȬT�/�q	m�0g~��g�z��&��=�E0�;G�^TM�y��!j�����+��u�f�n� �5M�F�N�.t-IC�̌�5ń)w��4o8�J�%$BiY�&��U�L6�N
�Xu2[�oB$�&GF������|[��a�/Q:��=� 
�`^G����0;���#]O9I
��Zԗ���P�?�U��7����w���0&''Q�v����\�0�v�H�a���wL\&�m(�K�5��ڹg��q��)��6���e%�B{���c2�[::���R�2�)8�f�>�a�_j���c��ٛ��l�[	1�?�,'�^�:�'�;��nR���ެo`���U�2���;z�]����=و[��R�P���m����(u��2���^�K�!D�6���Ez�����K�� A���QW���Nu�{�d��c�a�1}T���1��n�ʸ�E�D��l��w@�����0^T��/>�+�تƍ�aj7�r.!o��ۣ n���#�4��[�&b���gё�'��w�ܴ"�2�qk����	FH��wS \XRoo���ۍ��kq�'�>�e��G�o<�T ��,����vYa滋>�ׯy����h�&
@���$�����t=�a��JSB-��,�y�~@�_�ەD��|Az��x�e�nP#!�x���ԍ��O�ufA�Ɩ��p�*	�&畜6�N��i�Kj+���X�4���]�/>��o�M�xw���c痩&hX�����D�N7�l�G~f���2RFդ\�������:�ZY"
[KNҭ���§)o���"��M�/���@�Q0q��*��j�@x#�:F���B���X�t�H���_�W7-��HDF�10@� � �^%�=���'w%�D��\E�H=�`S��Y��~u1�;ܳ��t�	g��/E,n\�'
�^�6�Ab��`9V��&z���T]���v�Z.�g��G�|��q���Ty�:�i��*�-��f�G	����z��]|��8�
�w�M~چ��ۢ�S��ax~o�s ��#�)1
%��W��yu���vF�"k���b��F&��i������VmV����&��Q*�γ?g\�����y"���iˍ�l 鰰��<I #1� F�\�r7[:��+=5��%�E�)>������M�ZK�>��v��W�̼b�`jc�X�Q2�iߋQE��S�H�߾�a�3������z���՗f�_]g-Q�n �7f�ū�� ��M��DT� � <;��i&�
\��}ԭX7A3_��G��?ۀ+¹$�EHQk�%��L�kT��nB��9`A��c��'��7��Qؿhc����!�r�t
�8��Īy�� ��@8��<~�����/捒�j�#��6f��@�G�Y�%��4l0a�%�E@=+M����s#gI�B�[I�w�&�)�+�������[9�G!�-YU:_ŚwdP��C��T�
����y��'�z�>�Dě=���3S������C+���N0X+�Re��5yM8�d����+�4]]���z�f=0���x��̽���ϊ�~c�ӷt1o8��3�J�7�`iz]6K�C(��RjB�u��\@kߩp�<�"A�$��p�_VSBlX;E����a���o���� ��8�e;����ݕ��a��s'�B"�]�f�F��a��ܝZ�g�r���]�2"�.�RK�ɘ���&� r﷢�$\n\���p׷|KN����c#���%FY|���g|��@����#S]X���H�9븪��a�"��	�3�1��4��ɀ��z{��޷%Z���4���b:�PEϵ���aAy�X�w}K<$��A������R�;;sVXd�9�����>����8J]@�#9�-�^�Hr4|>���s�-�G�.>؊Dܳ����̱�z4��=P�Ǭ���q8s�Z��@�^���	j�F��~8d�4v��T���(ʯ��')�҂�~O�� 0���Yhw��/�Y�o�M��޴�Ąs�&X�ljF͎;�jvm�h�Gr�*:�o����E!�Q�ِn}:���%��O;wW��%�Q�
iי�c�&�s`Ȯ�n�����̫�&Ő��f�cii�A]e �v���nQj/_�6�2b���'�a�Sצ<�H��Q<C���;O:���p�mh���v���T���|M�����N쫞�}޸F�!��� D0�Y���7�ﭫgVU��ܥ�4��"j���,hj2sc�"���1����eQ�{�����Mi&���{��b��(kl� �zP	�d� �k�Y3�q�	�o,��N`�E
���1gy�2�?�!]��V� V�L�s�61�� z��80����0���:��7�D�cs{;��{{�,���� _~�Y+���?�����
�X{���w4��3��3��;}���Gh'��U1��@�-@ӗS�a��Z�^ޙ*7���u
����s������gt�uS[-}�����6��9	�^(Z�Qj�y��n�b�jfW>���p8Y��u�����L��ϵ���{��:���g	=��  ���=&�r��m����g�ǳ9#��$���}.�q�����8�d��ŸŬ�u����D�{��%����wHnH�������k��뵁��L{�����7�"�z���+��pu�C�dc�趄����£�$��A�!�I�~x�MӔ�ǉ�YK�Or���޹U��O�-k���:�ce�Q`���>`�
#��s�9g���,i���`x��簴�+��. �|�z�ǣ�O� ���� &���ݷZ3��	�>.$u �tgz���dg�m���sf���{�-��4��7�I�j�/�\��LUᛴ��ظ)���%�|:sMl�.�b==�����Tra"DڇL7���ۣ���bll|�gk8��r-`g��=��]e�:�����u�����iO�	���qjg}4Q{Y�̨tN�"}ǼT|Ǎ*�6��a�*
7�6�0j��E��d�q���c5�ќ��ȝt�����(�ܶ��	�!A�Iv��v�a9c/���(������n�(�&���b<2B\��^���=Ҍ��k������x� o����i @���$�� ��k ݤǮh�=8(����(�MN*��	��a�Y5��j�0uk��e��o(&�/rl�ȗ�x��/��Z�y'�g�.Rwdb!!�+�C!�γ�N�oH����1_�� p��/9~�Y��j��8N�����.�W�@c4ǻ+�N�m���`iCxǔ�n�{Ev�ۓ����� A����,�P-���x����Q�9�~�����\J=&a/����7ٺͦ�԰ %ſ�V@���Ҷr�l(_�M䨆R�=�~Ni���=��>�mYʚ8�s������2 dl5�N�4��/�r��)�P}c��C�����3�h�(����5��������4�x���pϿB����GJZ�j����%���/z�g�)z�Zs=SIy�	��[��s9e����2�Ł6P�+�ɦ�G:�|����{�s�_.:������?���=ʤ�P{�r\���h�Y��nre�������2,7��a�A#��K���xH�����Qg�݄�^a�#�Z|��֌5E�����A;F�H��wD�z+#�5B^�Χ�
���c��]��1��~����9�:e�CV�L[~�խF�aj�g��ck& ;Q��n�ӑի�Q�>�մ���2�O"�+��sX�<ｘjr��>��Jׄ�UX������\V���ˀ�]`���*����e�9H�0����?"��SHq,�ɧY��E>8_��z�'��]|����-]��K�H�h�'�0������<I�r���wԤ�glp�|w�pZ���ȧ��C��ݰ*Yi�n��<�i���E5S��L[?�Q����i;#�ϟ?];��d���𷷷�<��3����)��$��a��Ȧ��]-ф���U}Ҁ
[ۿ5�S9rp����z0�Y�Ko�!��ԬS{U�y����$�3"+Z�os�N`�A�$�ҷq�|w����L���Y��^踽AZk����\Tdd�ǆ6���W�X��w@q�/5s��Or�ij�&[UbU���N�SƖBW	m@7�|�Sl�)�����ᛊˤ�}���Y2�[�YrM�$kq�� }����l�x <F���>a�w�����; **���OR
��<F��z'�]��R�e��V��G�
Tb�r><���ZI���'22�*-9-R���k*㻴���hBm��I]��� Z��|z�<�@Xȹ�'�.
�/�jG�c���,Z��D�ƼW�-�H�.�wjYx�m8t5�Wx��b��f�@{mwAY^S� ��:�ah�^���i�ݢ��r>�Pi4 �)�c�khT"�\�q�����hGO�v��Kǅ`|����H��hn=�"��/	���"t�fڱ%�Q��|�9~̳ܵ�� ��8BxO/�b����[*d]��ŜkQ�񰴞�!4��ss�ewj4u��u���h��{Vwe�$�9�E�X���>�9���{�U�hC'�R�����q�����6������{â��}�.�P1a�ȳⰳV�x��Y�H�;���|L3�����y?�W h�'������nf�uML����Ff��p{����P����ř<��FV�C��ca'�&(����p�ɬ�s��7�ϑ�8�!�ok�LoKP򽿪q\Oz�C�:���t�@��?]Ƹn~|s�˻��i�Ա���.`I�z���	���]G\�|�8q�����B,r������Gu��B��15�dt�K�|@��Y޸�P�d�c���,�����VRڿM�a'�y��n go���>���(3}��A�-M��#� �k�!S��U��r)��R�\���ISi���%���Y��@(FY�rV\���1�$�ت��(��y��霢�����v5�#2��~��M�B�~�q���4�F�,��� �9�����'~�x'8�Q��:��sV���TJS��v�p�sUd;����޼R	؝N!�Z��G��*ρ57��u���Kž���C"�3m*�Wh-�H=������\J�Y署�"��3a�x�I�h8h�7Α%��p3����[��t � 9f1�ٔ!�g�vvܨ;3(©��f.�+M��~3غ���1񖸻{��j��|�%��NoG���M�b�c��%�?�9a�A;�PXaC��
��.�p�_�
B��M�Y�Q�1�-����AGIEK����r� l���&^����B`��05���.g8T��l����j�ȉa�?10��@~�q�x���C��5�Q���O�ݦ.IA�IȽ���|.����0ʷ����h��U��������	���gѮgי�Y���KB�W��[��&�]4Z��4����(�B��^��w�!XR��������p��n7y3��m`������IZ�OШM}XPc^Q�GHB2��]�i�^�3$fz�"�˟PK��a��[��e��ȕ�kԁqQ{'���`�Uy����h~\���G�!U�UV�$轴 P�{�T�>�ٟ#:a>��F��:,{�f.�|��l�a�L�g��z�F~0b���얆�8{h���q��L$F��22�������2G7~��,��:-E�vJ<:�s�C�>b���j��j����+������z��m��T!9��Ea`��7�yZ���DU~����o�Ht�������]�������"w-x���̺��ʶ[�� �ӌ5�\0���	��/!����_&"�q}(0�,5���_���	�q����H�����3���XX���ĺ�Ԏ�ʄ��S֔�;��A�3���>!��djEF��/���@�1�#�o�dZ�k��]g��p�[wh�ZJ�] l���^�P�E�9L�H�Ѻ�ސW�P���[3�^�s�������c�|���-���1���0��'蘮ʝ[׻b�>zm� h>�V^��a�J�^���:�s��[�įu�,�'e��f�a���9ˆ��q]�,i�M�@�8R!wn����l�ov�;��z��TX��A�
F$���3��T			� � ��c��1���j��T���ü�K������up���CJ~/)�V���(��/��)$����}PV��S��s�>a/���g�ȅp*��oj k!���/��w���j_�n+��=7ί��%m[L @�����k�v?�aK�=�����N�ؠ�����v+~�
�3kk��ʾxFiR\�љ����~�}:?#&xC4���%��
J49M���xƂ��U5��:�0��K�>�f�j���5P#Ǎ���!�<!�mt��C�̇z�U��K#7^^Y�Z3���\<<�&�gF��bmr|U��?k�=0 ��&ۋjXr���Guu�*���q�??Ҙ����wl���e#��*RL���C����0���h.6�0�����@4���[�h�02�g��"�X]g�Q ���l̘:q�&B έQ�_����/ӂߏ��j�	 +d��lw��
�߯��9�7���n��u��k�?:>Q��7�0'��:�u��$y*P����n����C����g��a�<!��4�a`�2ԮDW-�'���~���t�|��;@�Y �ִa[�����Yom:˘)+
F�S�90��e[���F��b�e�6d���@>�G�e�bW��;��4��`��a���̯� �0'�l9��/ĹJ<��fYf�w�!u��μ��
n��`�~��l[����ՌG�!-?`�Q�>?�;.:�$�+98��]���vQ�3��T�z߷.����N��OTSْ�'�mj�?��9[F����C/����!	g�����ub(l�70 !�����g�����cD���m1.)�cM�������JJ�.�Q,Z��li�#�Q2���ђ�>ƭE̮z�{����VG�f�����V��x�l����Ą.}�!��-����VsX�}4�W�w���5A��c���f��hGƇ��}5 {�<�yC�̀�9=�!�`:`��sKj51�8��l�~�h�=Z��xX� Cͮ�i� ���n�4x2��"��-nd�Y.F�S���e{���?j�\�B�c�E,Lt��X�0R�J�����.�!=�|�R�`���9��Ġ�1W�+e�"�\��ȏ+|ځU�����)%w6�i"��������{l�z����}Ԧ�$K'��qx������̣�cz��(&?�����g�֘���Y/����rI���g�f��Rj(".�z��%�s� 2*
P:/��@��=3����(@@�l%'|	\�n�@P�Ls�nK�z�yۭd�i����v��t�[|�橛x��n�v�wX� 	�TKu��4���v�..}��}n@VȒ��/z�&���Uv��Ӗ�EZ�`]L�t�]�P�>����Մ���w�H�4�$�!���Q��j��c�ȵ��R�9�B�2�����%*
*v�%*O�=M���b7��k�}�2�3d (���n�3��m���v�b`a����my{�d&-Dؑ�>3��91�!��Î^���?%1��ALgko߹���d��km-��Ty���N5�D��4>?KQ)-]�\�~��_el�~MϺ�1�� x�vBO0xem Y���!�:<.��X*�c~K8LW�4y�T����:+�;Z��Amو�MiRI��߆�k*yټ;��e�0�1R.|Y����[�p������Q�YU{�'��6�Oϔ���1r�����NGz-wF�l�;�:o��� ~�MQ����7����?ޔ�n���X�/ފ��NS��b f#;;{s{[QM�
���`���C:~Y�r��>�&힟&4B�Wq�Mu�-�˭��n|j
��R��!���h&%�k���~`+�e��n��]ޓ,�٘ʸ~J�!&�h��|{	򿻸�<ۀ�o�՜w�.#ro� ���rFF�M�{��7��y���vd~��|�����"����:�"⟹v��	Jt�����B\	��07_:���P���ca f��g~��'�G6��kj����<�����v����j��$v��s�I���@U뮯#�?:��CF�#S%�טO��������q�c�L�Mo,��V͏�V$���za��/9��
4�6�/z?w�Ċ�v���h�Y�2�O������,U55A99����";HB9�ϭ����2`�l�
�����Mc��%���y�w�okk��D��(9Z��Z*=##N(ţEv���?`JPv���'�f��-HʧO���sXo��]�z F ����T�уl2��Bw�3Z�����I=s�H�Є�����"��J������Q?�d���G�!�U�Ѫ��"���B��&9M__I
 �(= }��-�)�{����.ˉjL�&���{�(}��	H��&O���!VR\TQ��bi��g������R�^7߳�1|rX���uf���gxQ�8�-y�8���.�xF& #sX��z�Zp��t3R���n���ˆ�:*<0�h�@�{�V�\ ~���SB���&b�?�W��3�贐���Eǝ��M���n���9�1`�m���qt�n�3��'+]��y\�	<%��7?���z����*��@ش�Y��{��*"�15�o/���X����q=8�x�탨�ܖ��kd,?�1V;�Lw�P�X�V��%�}'DQ��v3��E���A�P '+k�f�@.�w�bo�m	����t�!��-�9�iq8tu�	L��8v������*�׃%Ա�v�^�w.>��k	>�PJj*
}Ξ!u������S��ӡ�m��^�13w+�(�
LJ4�>�	���������f�\>l�szv����//ޛUl"6
- �[�*v�U�i��z;���j}[z9��yʇ����d?�)dlL�z	G>����qſ�:��WZZ �8�iUE::I`Y��	Ø��R�A�旅��υj%���{^�@�7θ�w��:�8��#��oO�r6!�~?o��/���U7%,0��ծ@��ݓ����Ɗ����kh!����<-����`L-��
\d5}0<b"������NQcx+��� ��.��s�	��v�-�^�������R��}�z�ñ��Hb�gX�ueea�z��3ҁ�:�)��p�ߟ�k17x��#��l�M�3NW�d.�!�K��Ӈ�󀠛=�q�镯�����J���n}M�r�曱��:�h=�L��8K���`ߌM./�� �m{�\�,�c<��be�y�r�C��)&�Y�����ʼ��6����O��+6� �w���t6��Nϖ\V@�zѵ�R���p�
���= ]`�DH���6���Ug��t�-�*G�2����l	���|�[�m�7��y`�]�fl�=9��/�'����e�/aiD�eDǝ��M����<J�5�O���+����Q�d=���� �r�t�L��H�ï�ľgVY�|�c��D̥�l"��!��/ pn
��-HU��gԳ�~������8U"Q 2�׏��Fo���i����� ƭkcu��7��B� 2�+��g�QFei�����T�j�%�����4E���c�t�RV�������Ys��ÿ13�8���p��;�	�W���/�S\��R'�C&�����9�3�i�gg�Zb��2�#����2��)�T[[���N�f�/:�Ќ?�� ��b�����*��1�v�(��]����<
(��Su�B���ؿ�����]�����#[��Q+��?/��O�ڒ+tGe�!�y�0���gX��20y7�|hHNE�u��Vr�/2�&���n1I�K���F�g����"w�ܜN[�%r�K��vF���+9���+�����DC����w��=>�,����ʪ�k���q;�[�2^J�*A?|��S�����p��,>A3��o��IJ/C�;��D��ٟ#��@�.p$B�!���l�pש��t8���kM�]��a7y͠�����V''' we�:X�)��Q�n��2�Qds���.٤1f8<T�<�c���`�
]9��J6�##���o�.���lcNT|���&oGϞ0�z6	�]�*q#y[~�C�l�HD���}���DRNߧ���
��|������������
�nE��@�����U\��*��sL>V�q�^Q��B��s����4�غu+)E�x?œe
-�Y"J�}㦦�<���yï�܊bsL�Ē1�H䁜;��'nSؼ\�;���Dp�����{5����Q�����7*�N��Ɋ9�6�ea�m)K���Օt�pN�^�*m���P�0��'ŀ�j�NSJ1��}��1��y��
�a'��u���V8��{^G�^7�����P�ii����8�$�ɵ�9�[��h���s$5�A�"W>�g��?׸p�³خ�pq(���U��\D�I:=:�8N��?�z_&@ajk�]�B�q��|Kjii	H-^C���J`��\��ѿ��1���A���>��6��=&���n�����M{�j���\��A����.g�e3�I���/q���a��aq�7��Րϛ�/�#
���[h^�`9G��;���!	��s�gE�r�\/ (/S�j��5�,�����ߛA�}�$�z1�0))����
�4J�fB,���Y�?��&�d�E��<�ш���\���.y���`j���"�NU4G��
[4�tD<m�A%����QR��3�8���|��3Ab<s�:{������pZH�#�ٻ4�
%x��tȟ���3����o�(n����oPy�����e|H3�]TRwݣ���}WT�UW�����X��G���~����I��KX�)�#�I���{�}e��SF�����E�?��1M��^�1:�3텑���<}��9�/ƅ�yY��}�
<���o7�vE�!�A���5F҉���%N�K<bf��P���N�;0���*�wۘ�^S�.�妙4ʗ�.m��:<rt	��Jg�I���>��,�d������\%i_=��� ���4�y��3�����|���x/���h�-�I� !������S톁-@�GG �z���s��B^��u��z�;WgA�=io'�<	�k��ГAȑ�[�B30�3ꀩ2o��pIaFE�����壩�� !����0u|t'z��,���xM���"�|�)�����=*6�:&f�G��m�_�.g���H�n�m&��&�lV~�!������=%���s*"x��2��ߘ�+<����c���e������Y�rߏރlLDk�ࠋdu�#�F�.�x�vʽ|����A5���M[�4>=N6��@Q�� 韲a%Gg(�C�p�I}r3�q�^L�iǲHMH��m �{|O]��y&/nt����˜,]�'	��8��vj�����cofNf��%s�"��n����.=_usb�{�h����6G/�q�.����RzL��m�Qd糙u0,�(*=@�fZ=�k��v����^�s��>�'��#���d�Tj��<]��:����N3S��uŔ�/ßLv~[z�e�Y�T��^v����Է>�<�<���U������;���Q�{}�� q�!=i�jUp���������hh/�WG�|]_��`�J̚�C�o���ҒxQ��3��V`��C1P컑�	e(h��W��}t!K^rX7�U�&Q[*�->W�g�@D�&�{o.�������
�3j'�#��yqjm�g���SW	#:��Ej4���3X�=��w;kb����2�MJ�߭���}#�H}��iY4�bz�7:y�Iʰ��H���ёp���|lb�!4�q�[AnKwO�#A�V�
�<KJYF׋���Օ��@��ä���)����#d٬I��ԨA�jXtv1���L9�(�������O�c(w�6dF�+)�h�����u\7g�^.�)E��y�N�K�V���/<��Ǿ�W��(Qz�����;�(ʻ��8m2I�\(�<�:c~@8�w
r7���o+�_ׯ s�8�ҏg�O�u�4Üמ�z)�CR/����s�	��dk��a]�����+湳�܆�Y���$�h澩��4�ݬ8���nҜ��>=u!,��Bn#�3�s(�~t<4Y5�.^�uv"W(�cֻޅSآ�~���{����X� �eח`n����*\�É$PouP��c��?��n|����@����Q�.b��}���r���|��Q�����0����a��2���M3k��wE0V��G���	�b�lS���b��&���TI .Q9�������J0�Qw��&^�/C���Ĉg��",�� ���2W���`�U�>땻����,���%�����|}d��� ��?}�Je�)<R�R�Xt�0�x�)	��(e�^=��� �p?������-J|L��Q%F���?�'І��������'���E�����*h�s�]ٙ��� f=®�q�8j� =0w�[��ӨB��H�C}�	��љ��~���|%>�<��Q���������k�;���n�HiҤ)H���&�w%4A@�� 
R�&��� ��Ih�BI(A�=����˛�a�F��{�9�\�����ۿ��<K���ht.����"	QN�*��p��)�����՗R�ݽ�$}���/�u�f<�����c*4(��4�6@�`<##E�{08�Ϯ�$r�Y��Uc���;�l�'����%���_��^큳��v]��n���g�Y�>էy�O�lSW��u[i�S�zJ؍l����p�l���g�޻�8s&�[����ZP�U���>�񪕭�#;9[T��d�h��Q�#;���`���>zT�W������������o;d�
aI(��(�6����U#30׏اo)ޛ>��;8zfs��"�nf4[��Eӽ�!�^��M5!讷��.�e�h���6}d����� �+ܷ����%���炣�WXnP���gJZso���}������η�����=�rk�������7�,Jݤ�ކJ/���������b�nBk?�X���o��j���}�{E˭�� �`ŋ|��F�2�u<��ci�-A�t3��4^O�Pؘ�;N�u� fbW]�S�V��8�6��|����+_���wmxO�}�2���>#���Cj�0��F3ڗ�;lV���:{�����\��R��X���3�<�uc�nX�)}V�
P'��՟��C�ZGa�:���瀑ac�sw�p��k+Ò��	5 �`G��T���K�����w�]�6�~��1򼆌\A�f���:��׮���
{c*�3`w�t��EbG�]E>�׉nN>�~ȕT���	�_v�zz�j�>c�*��+��Uv�r���C=�8��mb����6��+�74S8f�M
˻0��o�����O�)����ɤ��9��9�� z�l�����J�a�������}����K��a���x�7����)i������Wb�+��"?�"WR�14�G/y��~�D���	�l�D��O�*�D�������f)��w>��
 ��N�~��nc,������$�\��$�R�
ѷm2 ��h����y�Ω����W2���z��-�/{SQ���V�+~v�bշ�d��\^2U��JR����(���\Q>���T��X3���1p���aER��d���x�8x�=��A��J�R*3�7˻�ք���<_PO�sMX����X8#u1��������P��OA����͡򟋧x�%�ºOw� �Lqɩ|�1/��wT�uG�ֻT<��>�z2K������-��z_�pڔ��I�)?�E�C���'W˰����%�y��m"0 ��hg�N2�6d0�X�uU����<���2`�6<����16�F$#1�l�#�;�lI�h��źS���K��K��Ffg��S�; ��u��`4��N8j�<�i��C^�-�O�X�M�n�OA�2�\��x�a��-��L��L��zqV�xH�x_ ��@��W�^��'j�����g�r�m�bً��eڞg��H�D>��ޝ]9�zB�(y�5_1�I� ��r#�~��O�#ۃ��������T��zߛN;�˳����4�����C��CNO��`Yœ�ĥJ�$B�3[��\{�g��\����zE����6F1`5��4,Ai`�_�+�':���p������e��1����ѷ2���X܂��'���J+j���Ey��{��U6p�B���t���y�~\�\<pށS·��" �w`LޙM_�
���X�CEa�òp�c�[�xk��UP�>��qv�N/;��O;�!�L;%0ڑQMC_���J쏨K���ʹsڻ_)�]�ԥ�N���+�J �*�0�(K����L��#5%���V��L�jn�bއ�[�#��s��Zʾ�ʹ#;h�߿"}~pɪ��PhO�wP��s�I��UOk��.����V�zaQ4�iַ�&�٠�2��Y��7h~K�m��G����W?�g̈\��y��-ғ���؜���/_EMkc9t�Hi.@�7����+(rܬ�`�(�Au��R=�,r��ҤxX[����͞=��7��S�}���4�Ō׾d����ټ�y��� �Q}Z��=#���U������O���oayQy���dۢ�[~�q�=<�{y�0[�S���7B��!ݦ1�IbQ���p�&Q�}�0�9)ЈBa��� g��v6;��0���.ϰU���o��'?�/�?Q�8M۵���b�� 84��P�AIz�tj��f2�y<x'$ȱ���$u������_�3]|����f�ѭN<��xl�|�s�Uty�}?+��Pp�(dS�ЋM����^Rq騏K`�5dag��h�����c[�לa�Ls`�P�-��Ԯ���3r�@8�B���9����a���/�%�<aS�{'����P-�?�)(�L�)���̦��@+����g�	x�����T@n8m�����k���ƢΉ����:��&~�GA�KCd}ξ�i�{%T���e(EN�,z��}���&O߭J�?��O�4b,�������������7��p\�mmgƥ�s;����\�^���0�.`��z�x����_>oA��n`n.�t���y+l�kv�萫?+߼o��q��?�G��ƭ�GA�A��g�r&��?tƋ{��T%����߈)�ٮ�_L٨٠��Wy/�y��}�pPab%L!�Q��/U�n	f�}�5�q䟻��x�+�<�q;l b���`n��v��E�b⻏��t|b"���j�Lup֋>�s�N�Y�nЯ��i�.pL/�r�B6����2��@�c���.��E���,���������w.���z�{�,�Cҁ�FG�mUb%�O;>��kb �O��犹�`��BS�k���k�Q>�޲��9�j� �߶~�Ŕa������ƃ:U9=cɤ@uѤ�/�/k�����BHݵ���#TFs����=��������/�Bq���ӎ����Kh��/#b�����F��ſ��]ئ���}����uf���%�˄�i���n���-�'�(�R���7��NO�e���b��rZ�	��[=~�_�I ���Z�QWx��ٳ�z=��|넘��R�t��4d%gw�"> �ʹ@�9�+"�z�C��7�@�ˉ�*ǀ��WTQ��Z���ѯ��5��zZ2�E7��[�}����-U;��'D�&hd�KL�˳[2q���1��|B��0�|���#�Ώ�2��JG�r[^;�怡���S�ҕ�#}R3�q�	��Z��ª����n���ɍ��d�PV��t����6:��z�d�m=�%���y3��X
��z�P/��51Y���b\||�p��P�$��
�j��7��^^c{�u��u�ן�U��d����yDC�#?B��X�8���!y�L��$�ρ���s�3x�d����?}=Uz�,P�\��#
'���fl�ή[���{��޴T�O5�sr�@y�;!�����s���@O~U��� �8���{���=/�H�RÈ����8���IYe_�aT��cFe��T��ߊ��A��~X�����#�*��).�c��JFl���2O�\m�ؼ1}☦�t�~$+����8m��?/J���1�%�p1�Q�E�Y��~�Hv�L��囓������p������ʃ�[*�5
�Ъ����pO�������Á�K���>����o�
i��覉UO�3ԸH�_[s"�D���wqw�tM/��鷃, o���@ؽ��XZ3�A�U(v�y-�n�pTOg�U�����o����w;���jE@�!��U���#!?o[R���m���W���^
+�*VQ�H*���T�zl�����R�Q'��nE�(�ϩv���>������<�	y��Q���r��pta1�?/K��j/d�]��S����YzF���ě�ra&҅�5����8G
�׮���خ��>k|�;,�u�u3Smm��)�:C��7�fX��Eg�.�4`r�<-9�~�L0�my�z&����K�M	�n��&�#��G�Zp[.`�ڌ��|��2����_�Ug�/:}/d20� �i�P�M��"�$O��(~��
�~|/,$���"l����6Jm���!�X�Y��^ ����]\]��������{�	[卍���*�~�~�2�u�J�ejZ� 6���JPȲ�s�r�]*�3+�J=�q�ڎ�0�K�Yuh'~�F^��}Fɪ8^)
^��o�a�^U��;|`��6�������V����:|;F�v�
�V���z��a�i��P�v���fc�*eea�'�@�ח���O�?�pO�~v/@���K�;~T9	{~^��NLL��Ɩj)���j�h�%=��U��𐰅�9��b�g{��Y�:D2��
9�~a��k	��p�X���g��+��oVɴ�=0��qP.E�ĥ�l�%v+��_Y����������j�=��;����6|������"
��\��o߮�>ZDJ�Vb)���p\)>`����d�r���CӢ������]�t������s��y1�'����Os�ӵ�m%F�!�}⯿2�6a�up���Q�:�Ϊ:M�f�iI�d;��lX%%�-ۄ�F�(��?��{�/J����b$A��Wb��@��E�fHx���eѫ��Z���U��B�ߓXo�e���V,)�d���q�G�����2�fdʚ�"R�HǶ*��x"�%N3*���>  A����}R2�0��~��Ù��s�r񻘬�N��2z5�t�ׄ�'i����N�Ҡ�SWS�>@��φ�_�5�	{"��E��b"�i|�Mu�`�C|����s�W��O�j�	�q��ƭ�ǀ��#�w�)�r�F���)���-���k�X����Ё\�O .&;�]a�^��3f�#x/�7.�<��0x��e���2Z�х��b��.�Q�K���XWOT�9]4�JI�����U�$u�#n`���w`j���y�vx5+��ߴ���(Q�"Rc��ܐ���Ί�=�\z�&�J���6K� �f���1�斣<��W���;�A	�>�p���*qCr��IP�6c�u�fլ����ũP=(��я�{�7�QQdȌ�Tcܕ}��~���85���Fأ����	�f=���$�H�-������n�Z��!�C�����{�|QO]����/�H�����ϾT�_d���-	�=���q@>r��m2�e�Ѹ>�JSx�mKES|'�HM>������)����g���`��-f���:tD�_lCq����1�эzP�@��gkgl#������
ߪ�/���b0�uj�����H�C᫸+Z���o: iJ9���HʓjF��DR���Oڻ��hC�\U�g��$��s�H+�\+��j�I�[���>�]8t�]��_2n��X���,:��-Y,�_�r���1�C���r��{G/+�u�p���O$7�����&%r���;��&�~��/E�\E�F���y��Y�t������lve�z��k��"^�zT�5_��N�xXW�ib��]�H1p���|�s`�O��1�-�Xxs���8܂�Ȍ��O�Zƍ��5�J:"\���ߤMW�.H1Wq*�cp$eV�U�+Eè�T�os��h����eq����O�fm����s��M�2��������d҅u�gjs�T���t���{�����m2�J[�	9*+�s#��F�,���b<L��CQvC�J�k E��le���۠�m��T�<��:ܨڶ�g�a�ߣ����< ���L���D�}z���������#6�S+[ނ�� ��Z��Na�9�����vp�\*[]L�A�6�BD�^���Qўch1��t}����\&���5a�od�9�G�'&T��Î<G�e�@_��&*B��n�
s�z�.��n~�Ӓ?�1F�q����-p74�n���:3�mz�#��[g�?h�b��\�$l�*q����¹�����ء&A��$�iE)u�����k�7Nῆ{�Eu*sf���F�iO!<Dd\�Y�$��P��n!d�u�WkI+rtl�㠄���������Ϳ�39���c��=�þ��\��	�l��]x=���-ʑ��
W�,;��Y|zRx�sy�;6tug,�p����k��~rT�>L�i�� G}��S2��3�C�Z�}��*B^o�糮3�>��/1�x�c��c�C=����$�� >rJ���|��B�y��ؓe���6��6��D�?{>�<��`I�ٙ8?%˟��ė�/rT�i�r�BG����*�q��2N��;[�a�߈V����̓�k+��1Qy��_�	�ȥ# �räʖ$+�2"{�7�bE�*�����k<��f~_�8
;E��v��5�^.H��t&P�i��\�Ou��ؓޔ����Y��lz˺��a��`c���.,��SK{c!R(��뒸.m�����D����s;���I�$2��e�Ӡ�úӘ��V�m�#.Ц�7`� �E�����>"�a�pP��#BPb!	�:}~��"�r4��*�ĉ To�ՙ�h�hrD`��MJ!'����5a�p9����sKTX���>;�ep�FϮ�1mt»#ۊ��5�5�25���m�Q�#W�b ����lo�?�ܶW@5�� �O�٩���|o_�&��^T�2���dU&��r��.|�%<h9��'͂��IV��f���z`�`9��&�l�ÝꙌ�f��&���i#�Ĥ�횓3�v�}&P��u@7����"��(��.����O`n�N�[�u���Į����0�1���!-.oN�D�Iw�s����gҊ7'}h�^�=�V&�F�[�u�~�_�|��@e-3�0�(x��]ce����P9w><����8�Y�����nt�����,b+�Q�8OgeB��������3��aZ+��=C�R�zۻ���b�>A$��c����#�O-�ñ�p�\S��u̅4o	�~mִџ���G%o��'hC��)�p���`X{H@9�k�D��������!�/��[9��(���Ї�z��`޽ۣN*!�磯���0�i^��#��p�(���W�_�U�}�l����u7�+�0����wu �7Y:��C�[' nA��pWݱ�2rpڗdr�o��!��6e#  �Z��z/��{��)�{�j��p�'���~�;�ၮ��;����b7�D����1��=ٞ(�P9�P#�\���J���5��_P�q��ν2%�1��+Po������0�x�	m��z�I*=
����3��7�y�I�|Q����X���ν6�D��)�uI-B�A�fu9s;GnIs�C':X'��@G�z#�E�ŻQ9f�j��&-#��LR�8�y
��2�j��I��#��4% T�nG'az�O}~�@�����GO���-�`��3Vv�磗��'��[��bʑ,e�Q[�A�3V�Nv���}���(�!�_	KоF�q@p��ȼ�S��m�%2LeK�������9������s�m�����M�|��(p�NG9~�[�dI�����4���3���#G@x��1����������4޵���C]�x����Ɠ��!Q!����$J$?VB�]��'D�j��;~'�xa2܇���бpQ:E�#��J;�����ȼuʙ	2��~Z���ݓ��̱��5��cIp�PNп��v29��o;���p�_l;(�LC�b���#� H�Z�ke�=Ѩ� �~ӿ3i��a�p�1�sӭg���=4�O���e�~:��ީE�������W�rX�G��|/�,gi��G^�[���H�3u;4���>�q���	�	�J��|���j�:��e
Yawm_&6�ǂ��u�����kD׹��G�\���`��eF#۲���J1��FG��/��v��.v�	��z��H�_�b��_���T~X��e�����*��&� ��m��[Q�4RG=�ܾ^?/P�l*p^���A�v�J�~�߅��^+|��[h?^'$�SJG(*3�k0�K��_�������󌽆b���XU�`�VL��%"����G�
`s���f�>.,(���sO���҄$ �`�b���S3�Yn!t{�|��dUs7_Ʒ]��Z�R)�r�np6f�&���*�&"31��f� �����#�\C���R�� t�@L[k�:Z�l���:����fΘ�	=O�Xr/�&�vE�����/nG(������
����e�����9�æ�٥���e_9��Kpŷ����w\�*t��_��"��e�[��N�1���h�//�.�O3�!���=�݇x.���儜L�H����[v���.�a�y�����G�'c �j�3G�t���r®7�3R]�P+�m�ܰ�����8�@��Zt���i��o=,O8��҆mZI��Uo����$�����:��|�\.;߀�(�@-��"����Կ�Л���Ϧ��Q:����ޏ�P�C����m�5�I�`ۑy���`հ���w5�Z~ƍBӇ�<j����]	G�Z�cD e���3�eb��=(���F��zj�"���w�&pI
�J-���[�q6oi"��U�`�i��ӱՇ��FB�K���Zܜs�Iћsc���U�`��'D H	�kΎ�$�i��#�$��B�4��=OT�
$��a,���i_���JVxh���'�������=�����IT��\57N��
D@��=�#�Q�UU�v׎�?V�.33�i}��gC�������n��q�?��a�qj���I��#�b�ښ�X�[UT�A�Xd���`����-�~��O��$�Zb|��9(\�p���s�16�����4�{X�g�я����D�%pe��,���w�;�K��H뢁?PBNB�Ph��y�+�޲Ӄ`�-�B��r���M�+c�Sr��N3���EK�!>�}}"�l q �+N�sJ_O釳��Q×��
^�DP���p+.���)k�HHO��!j?�IvUC�K8�t߿
�v�M����#:�}	�?�@q�3��9�[����֙@�!�U�r~>Ȓ%��'��G��FK��出�:�E��g�a�.�m�p(B���z3�U\ѹ*g�0ɛ crT��׈���G�$8O^���T���>9	��pa9�j�<��'�`s\�|���)�Nߓ/GO)e��L)����1A�h�h�S��fbv��5���0'|��ݔ�"U?s5�=L����}r�a�}A���S�v�H{F�Q��ř��O�"$�,[Sx���������]��JK�k����d9�p�h(��fn��A��Ĭ��0��⢜��-f��d]ϒъ�&��@�s� �����U��
�p"
8Ucg$��@�j<�	�&�Ɔwn���Fjp�5ֺ��s*҂�@/�_˃@̏�Ӷ���	���5��8�?w��|�z��.-�:�d7<��Mϙ������C�F��(��ef"��	)�$����e�Bh:�?��c�l�B[F&�
	�mW�2Q�|��[_>��-m�]�)Z�8W��z����yu_�84~:�d��T�� {������4Z�%@�D��x���>P_����J��D�V��c��3�@�W�n�S~T���6	�o�|`�x�/�0�GRo�ձH�q��?\�"n1䝜�_��g�9�;���@�I��� h.C�3�|�!b����&�������m�$B����>k-@��V��n)l�u�����^'*$Z���Z����a*-j�޶�([gM�3-	R ��bB�L�I�lB-<�m_0A~�.�P��!�(���~�gfˏ�7��n��j��?��Nd�'�*&��A'���DpC2���,�/s�a�v<a/�WmNhϗf�*C�0F;���O�`"?��9s��.%)Y�yX��x�5�r�����!A껻�����Lo�j���(	 ��v-�����dL�F�^�rjO}�;&����j{3�z������Qh�=i��*���f|@��$q�]�/�L:^��F�k��i��=���>���U�P�)>���9vi�>���Tbz���R/�`s�Oq0#cnۣ�!鿇�6��OWk�휂C9��*���Rw ��7��6g]Ź�9P*���C��$�_�T����ɒP��ż=��wͷfB��y�����!�/��yd�6�� G8� H�:��lM�~���=a.�4��@C��_�m���N/;��%�w����aa�ax��������q���0�)�"
_�g��G*�&9-8:�]%��-��A��?��n�=����0�8��S� &V��]�TZ8�la�=}���}���X|�$ՑK>��6v���_���3��]V�ҝ�n���F@�7o��;}΃�]��M�-T����?/����T����n�Yo%Z.X�O����Z2gcj���i�A�q;T �J��� ���Z�C�&<ƼkTG�K>��g�>%mO�ʏ���0Ki�2_�^�2t2� D�a&r���ڞ�R���Gf�s�4�H}c��"�6�=ˡ�Bc�j�L�� ��V���3���^���_?����!/O�`��M��,+A�PU���2����ȏK�Y��~�[�/��sU�o�U���K@6k9̟$G���9Z�ԓN�j���.���ٺdDwW�xS�@:�д̍0m�4��/������\�|P�k�C�,����uo�呿�P"-P2��"����$1��G�倦;���*�iH�pzjF �3W���3���7Y�#K������i�lOЀ@Fd������|��]����v/VC)6hY���I<57������mqㄞ({9��tPn���u�������V@��r���=uG2e�_�u ���=��E�*�K���!V���ݽ���]j��^|DC���\����O��+.��t�"���u�?�����mxK�v��!卂�Hh���C�����_K����7�=6^�ݿSU;��� |6�\k�;�Qfx�_Տ*��z��;���Jh�<'�
G��ٕ	.�Klβ\�c����iw���Rr9�ٓ��1��lA�B�6�b��+S�j�B�eS^��/|�X>τ�>�9��+��5��y���l��$J�էy�\Ϩ�9%�
�n�gA������>-�7(��Y�b���W6x�+|��O.J���
�j#^���"��o�L��f0����|��q�"��vK�F4\ѻm�م�ﭤ���:�g*���*�&LpM�M��t������Q+AҲ8�%��lm��Z!��V�b���>����*��&/���T�'���'y�>�ܩ����gg܍rp�W�M��f��hh*�8O)��]�:n'bg��WٲJ5&��±�)s�N��oy���X�p�
E={��6��kȖt������O�F�R��M�hm�_O.�
8��{˦���Y�OG�d�F�vnxa��˧���/����8��={DP�u�eC	�Z�������i��!%��ϪG�(n_T!�V߽H�i���*з�zs�[P6G*T����HH����1`c,F�k�a�F<���!r�]���ӆ=���[����!���@�����h�:p� ��=��3=4ؒ�ɯ���R^��=�}�]���?�|�{矘��|fa��#���cÌV��`�� ��|,PT>���y���r�/�fɲ���0�"v@LH����Q��/�厢ðS����l�K���B���r�� �D�}:�v�a�r�v�L*؅�J�����:m�������h�2p8��p�Ds$˕=�ƌ�!\w�z]d|Ѵ���Y�5��i!!	�e/L���:��g(,E�y뜬�ւM��8`݊��e��3��G��	5�3S��m��礐����-Q��H^h0}�L�_��cC�H�U!(�Pr$��K~���]6��Rn��-2u&\~�$ܾxثU?-�]/؃c�OK���^`4� <�K��(LP�V��;�� �~�ރy����Q�.�N�C0Иh~�����D(�u�Ҍ�U���:�$�}���D��~��Sh����J:ˢX��(���-4s]"K��A�⎃�����m�����b������>����Jr�P;V�$JQnA��wjo�@��tGBWiCM���e΍" 1����i9�Ƥ.����od4_�P���&������>�'De�Q/Կ�8��d�� <�Huc�n0hEFu^Yh�c����!��Vzbp~��1���ُC8O��Ƿd�MV�f����뻻w�k��kȏ��@ �;/ ��lY�_4�$K�I��V>>�k��1�\��ɟGv��q�y���fO�Iq��Kub�l+e��C�P�,��\Cj�˭N��K�����,z���m0�� P8���M�c��ٙ�C��⺡���,6���E�Z�	�z�3�N��3�oU��X��f��v 5��t0��O�a=����EJ�ƨ�[js}��E�ٌ��8b����p���)"��It��L���*ɭT��yw��ن�1_VQ�el�+#���.n�6��L�E�y���H�^���2��#de��CѡRI9HfB��Ԁ���į��E�{Q���P�b_j'�t�y�7z9���$o{�n�e�	��V�rO�I�ݓ5�SůS@j
?u�@���{4�5S�#�-�W	�ک���mIHhU���}C�s o��z�ߍtF���y2�:��/�D��f-�c+�A�m���{�g��H�~�m'/��_���L�����9���JH�R��y�}���5�~ ����(�>ʖ�وݷ1%���� �y���" �1 c��?xY\���&�mk�c�l��2��0��1��*Ztt`�*K�E��[�O64Ft�#{� ÿ,1�5��;T�ǟA���	�j[D��F୭�gZ�^m<(���6��OY�#��&~�z<3��B����+���lWIp��p��CR�ukX���HC�L@F������8���F�n��.ش�!K��kļ��*>!DUW8Z���of���̹;�����(�`�
O��>�Ͻ�WhP������F�<tJ,e�龰]=����$E
L� �����U��aJ��㉖mMS?�o�ً��-�vn��U:߾W�	�.��:QpHk�̘+��#�׸�`=ق�.�L�P���<p2{��Y�S����QlL[�B5螎��t��X�M�ٵ�tѣ��p�S=�i�����?��f��<�Suo��"$7psX����H(��L(�&_k�C�[݊��q�k�Z"��n���_El�\�����-R��~�Z_�ңs���5.�rYL���i���5���o%*����]CfRt`�m�^�\�ㅟ�<���n�R	}ڭxߝ���5����?e
�S����"�%��I���a�d��ѣ�Ͳ�����*��Y�'��/�HJZ$���S��(�F�s��?{K{��
<շ���x��x)�5��һN��E��ٿc�r�=������tY�����ڬd�K���UZ��٨3ӕ5"US���cC��b��U�j����7�*C��_W�4D�￧B��d��6��O�=+�ƶ�.�Yy��H�	)��q[;�>&c��66Iy�w�ꋬ+v`�kj��L��&r��VX�U"/���m�ʜ�9��I��
�U�:2��	+��*G��Lo�a�5��U� !�L�w�(����k/�� "*$a5��z���C��?=m�7����S���H0�����iS
�2\��F$>:��	iU��a�6��ѩg�5Q�p�d�����"����u!���
�N�-O���7L�kS��`hf��}���^�QآNF�j���)/����iw��П�y>�9[)0 � ���?������)�%e
����84����x�a��~���y�CH�8���a�����!�c�߿taD�=�Z��qB��sC�
F����d��E~��?�����|�[���A�{s<YJ�F��v����5�_���D>��-�'@�j��m�����	����?�a���q�!t�<�����I��Wm��,�`����͓����fR�Zz��f�Kt�ɣ���픪6�=��A�b���7�>�o{o ~�����$�t�$�y\D^IC���-3(�\g��m�i[�N�0���2��m .��y�����́�|ڣ8څ�y�ZTIY���`	者��`c,�&,[�#�{줡Η����k?�B4Qh$��"D6ꃩ����|�o�@��V��h�:�y���uO�#��q��RS�$lf�I���㞔�R�YT�����X�y����u�fpy���0��0�$��=�2�>��W
�z�F���*�֍t���&X�,q�Ϛy��	/re�(E������U��6ݭS���╅��W�>����YTgnh~�!]��GR����˹Ļ��vv��Ҝ�����Ø��p/��2��-P"�'^�ί�	f%�6
A�A�<�`Vb��ҀB������,�I���b�����^���U�(��C��8����o�e8��4��2un�ˊpKa��.�5��h���B
���O��\�QL�v�o��Kp��I�M7?HU}b
�_?a.f�u/|�w�b��xr��E��Ժ��EX`Њ����d���~V�(�_[pzKݠ�)��T�`�E��-nO�Y�咦ؖ\�'T�+�1�9����,9!��b����	�C��	R�j~%6��>=g�@KBW j'���P�k�Ï�\%d��ǹuOjP^d�qXM�ڹ~/�b�lY�&�c��sDs�%/������i- �Ì�6�c��G���M�I��Ւ>ߝ|:ٺL�d��Kn���t�"�<{��b�镐��;m�5�z�Ny��iN�iBrS���Qwr7�oT۸VͰ3��:��TO���X!���nݵ�t���F?�9t�蚤��I���4���	�:�Sba�����������)/	���lZ�����e�Ƙ�Y�2�0��R�JqD)�i�;m�=��f���2)A�W�v�����һg�T����M�ͧ�nd`�ϱ�	S\q��IG��I�x��j�Z���z�e��rf��)�-������0k�-������[;3C�������=���I^q����^�lҵ� �!����i2��(dў������4 (H�_a �v��5:BY��e�BX�Z�ZS4��D<)�cx�Vz�x�T��}3m�t狤��]wHj��[i��m����L����6����'�͸��"-Vc��c��(���, �Y�,��p޾4u�v�@	**��i5N=ywK<>�����q����E�hm�c)�e&�����̇)[ˆ(�iZY*��,��)QX�l���Y�O?0�p��	rݕ�{Dx�^�%��G%�?��{����=�����}�_����YXNy��j�A�z�媶�PK   J�X��� �@ /   images/3e1f5452-c6ea-49ae-85fb-ddf6f8b38dad.png캉7�o�>N*z��dI�"$[a��5d;ɒ}g0�RHv�N�l�ɾ�(۔=�a,��F���5}?����;����x���<�}_�u]�3����:�<�100�ij<1``85��p:��4��G��r������b�}�K�̗���;������xx�響������ǁ�H8{����z9Hx���&)�00\c�|��(0�0�e��]�ǭ��q��|���%���;�����1?���r3�kV�J���+�[59Zs��JiFt�Զ.��j������2�Xӛ�ћ�����w�}���HmT����ǐ|(�xz�`a��<õK��S�Gz��)Ji�S�F��"�a&���0*$���������5��٫��U_�(10l~||��~�����{�s3���v��=������_>�S�G='B>^��ݒ��w�����5����U��.g�8^I���⊻gNc�2&cK��˯i�������g
����L�}w,����N1���I��̢��,j�&~X��i���Lܒ�3n�����f�vێ�+��a𣾃��",'��L���	���f��q-s8��I�R�g�))j,*�8�3��E�l,�������(b�,1��,�@i�Zw������S+��o���(ySh�]xj%zA�ּn����NZѩڗT;@� ���FoW��j��)3�4���u��ᆿ�30;,ɨȖw��'�irj_v�����=#$�_�yY���c�KB\_���=Ζ�A/���QG˸l��~:��`���������D3���C�"F163��e��b�<��L��wsŗ����k&%z�F�7,�1Ț��M��<���Gţ��%4'����nO����e-̼;zS��^�e�)��h��Na\���Ք�S��L���޸u��p��J��q��z��;�:f�(=��l�ݬ�Ѭ�����̵�GWo�^�j��JV�[��	��lFLE���fy٢cZ /�d������&Ţ�f�(m����{�TJ�Z�R,�J���Z����ѧfV)Rv)|��tQ3i��!�u�rO�<p�����&�}"�Ly�_V4JV����;�ɓLh,/�Y5�CpI_�03 ���v�U���:�U
�/0���l5��=-.���4��M)��ؖ��g����f��A����8Xke��Ů2���!"����E��h��^��%WeXqe��fXTV��ϰ�����8|I��AbD�ʦ5��ӖIlR�ϯ(����E;��\/J~�?���Ye/K�G�S�+��]����e>[�i��SۉkH���#�legh��������hb�rZgwɁ�&��C���b�<WT|�;�K|˕�_8.Y�G��İ�ጨ�dG��uLh�z�hnoF��(9�7�UH�)������y?���՗~������q��=ӟO�h������8)!.���҅}�Z�����n�����m�>$%|nr�=��e^�5w'�\e\r���F��ȍ�$�N�J��l������3�W �#�53����u��ty�<#JW�&�k�h*}���	�=��Hhf��om#&�i�
�f�k88?���&��5������D�\]@���!k��H����q���n��\(���%�+�w��F�=�������[GaN��.�Clb7�GF����jE�+�`5�Z�\���}H�u*{+�V���
�OD� ntC�O�N�Z��س�g2���K�JX���\�P�7+���`�R�a���?����$�!��٤���S���������������1��c�#jX`ʮ��ʬ{%�ʭ��J��p�ŦJ��� +�ߕ ��RM��S��end�;T>{�g\�N�a&����Th_�a{a>F�Η�ZyDo�So������\śB��ˣ����oֲ
Y��}����F/��[��>��8¹P/sg���7*/Ǜ���c��EͰ���/��1���v��I���;�M��A3>s,��<����a���.2�L�!�ȰI�k0�ތD�_��*A�;�6�u��,]�]cV�R R��/�'ϋ��
��'&�/5�m��Zv�p�i��4|���.a��ʲi&N怣����*�T3΃xQi�4����1xܺOR��{?�q��5��Ħ�94�,n�l�� ,k�Y�+�,���]i�vN���v�O�:PֳW`����ZQ< {���K&�ُ��q"T��`q�������6�L�is[J��OBG��h�5[��M6�8k�A.��Ox��>EB�n�fl��I���'m#@���+iM�U!���+6c�S�x� �����w)��PܗBv�*C��)�Z��Ҋ.n�y'�/���P��;�EO��}<��
��?	���d�Ro����~[�,�Bxk�#4xv/�S8>3][#��sc���Բ�ٖ�&5�j/&O������~y��J�"e7Ai�����}�%|����J��(�ALᠥ�d�O��Ǝb�����������̇��ɓ������b���f6ً�<r�|����l����r�=#�g^	g��Ct��r7��e�N��)��(%(�����y�D�-c�{�g�ܾ����U�����vPן#S�F�8�2�o@E�쾼K�X�����%ԙ�qLOc����/�Gb�.l�T">I�|_�ո]�}[��&�mx�^�rw����c��濞-�����n�"�<���F����;�.d����_��x��d>�$�1�/�b*�%�Kj��L�	MG�4/�7#�C�� �=T0u:y5Wm�,�y�i��8k��,j��[�NP�&x�R�M	ր'��¥O&�����-��_XOt���/)��^S%Z:-�pO^Av8�pL��ר\d���'��h���7'�g��[i?+}�tdw)�5T�ԥE�W�nD��~��{1�oi�࿫c�{�ڪ�~�pW�UF�+@���g��Đ�p�� �G�Ċ���H�&h�aLϮ�[?�0�U��f�j[&�|c����6�u����� ��v�Ȯoz���Y���'��j
#=S���f��lTK5��y'�a�]���s����u�����!qB!��O�*�sG$��oS�c��7�VS|DOݷp��/�nJG9Ű=J[�T"�+Zn�s0�Tr��~E��z�[�ʺ)�1���룜��U?,�c2Z�ʤQ&]m�X}��=#CD��"4@�썂�Cɀ�J�a/'��x* ���^�HaĺKh���e�g6��6����~ɺ���i�ԃ��|��-Ō�%��U q����kFڰ����>%�42ڀ�^�����H�s�t��$rQ�+�2y[�]�S��7ɰ���ށ�^�W�ǰ/%�F,�)@&Y��w�Tz��0��ųu�)��O��}�G������{Ǘ\���-�>��=E�x������D�q��l��O���kJ����]Dý)���BV���i�����w�b7�0�rr�M����U���-{$��z�ےW��)��C҉2�{�0�6�����3ow��le� :Im0�X��ٛL�1L�.���v����t�@9i�����Q��X;��>�'�{�g5'�7���O���Յ�L��C��>VS'�#��⼲0���:�hr�F��=���h"w(�G!z�@mpr�〤�ZM��g���������g�Ceq��'����B@O���]�j�I&]�!��#��6�9���pҵ�������.�9g�u��B���)69���I�Z�Ԓ	�f�gl%���Ӂ� b3K3ź�=�_��({���L!Uh2�+p����>Q��ldA8�>ڰ!4ɅDz�]�^�-_����-����l��?r����ab��=1�&�9�Z�;��4)�Vg��7��~( j��~�3%�:���+L8�� ua�����A��d�ul6�2pl�j�>��<�=�ų��3oT��[�_�_x�����8�?!���${��-�g��p�⭴-�*�qMST���pE����~������5$L*[�\�9����6Ec�b~"�v6]��l�]a�HG6L�V�A x5Oh|~Ǖ�iޓulty�*z��Ku2$������m����e����iG@��P��%�PM6'KBF�����X=;�c��}W���y�}5g��O���|�]!(�	��[���dH�J�	*��g���T(-��)��.K����>Æ�l\��128I��5��,^҃����h6�V� 3w����%n����~܃R���^�7��t/�."�9���#��Al�Ffi]�w V<T'�c�V�=p�8���$�Xm��H({�o�����/*9�	[��Q��-�G������Tqڍ�4{���^���~��0S��b��H�$Q5���R��e#S��ؓ�l�e,d��2��As5����~��Ͳ:/��sj�]�V��p���$v+�t�-dJ�y�|��T@z"�>��rL8�U"��e<��m�;��3���l���}�]9��6��	��NFݣ��z�^�Rl>'�_����Z��h�hFY�f`p�@���V9|�h��X�%���dP�1AP~�S"�ZWe��!l�wC0�إ8�Q�a���v��ru��H�T�n��"�������zLg��.��'3ۆ\5^5�b��%�`��ǖס�'�X������33�$s�6K6�7��@���n6�����7q�wZ��`.�+��}��#@ݮ��M�i㵫��a�{�6O�=ԍ�����}pn,ٞb����U�.r%1t�䋙2\F�i�5��wWp٩�%���h�U�N�fH�o��(� �J���|�w��N�y�k��ӻ�b�.,����L������{#ze?�l��<�R�)Co�J�&�-�jq�+���[��IV���C|c.�RD}�+���{HM�8�>QS�Թ'����|�ߺi���,� d�t�_��ܹ�qfߩ_y��"_��wM
[9��/�N��4�����oP���Qe���'���/b��U����h�\��W �/�+�q�J?q(�6 �_�ݥ?�"@O_�TbPK������ϟ�lJ���y~�Z�uӬ]�3ό��P֍��/Y��+�|�f`x�/����K��]Y���6g}l8�z����A=�����o����~*;cni2"O-�e����s1R�A')�E��+�\�����^��CN3�����7�nW�z^�By��/�����|�?;����3�H,��f��7�c7�]���h�[џ�.Z��L{�b+X��N�����`w�W���z�KH{�=?�ީ�����D�N=��h�r�l�%�-]��xT�kD"�т(���P\6c��C�,�W,W�@��m��.���A��H�������x����{�AkX�*EWDx�\q�Ő�M��#{���V��N��u�H/���#'�Td��r���.��ZQf{��5C�?������&�|83
�(ݢ9�j���.M-�ڦ"W����>v��f����:Q�3�ݤ���Ț��#�~K�����]
�)��Fěc����P�9�����E>��1��͜�ƽ�Zހ�+S`�z6���B���æ���M��=�s%����>ݰ���6�4E�汁�)Gە�v�r0*����G`��o\aN���������B?����_ ����H�6o<�PULFi�!0�5�̔}��U}�z�;����?�<VUo��T�%j�p(�K��9(�U]�5Ė��>-M3~�q��!���xʭJusǫ�L�,zi�����,t�Z}m��P�O��6%�
��J�yT��2�ͱ�=���oTP��5�5Y�����\'�~I�>�d`��N�8��2�A/�7Z��� c?�?�z4P:�xɝ�x��츰�l�,�d�+��Tpɩh�1���h�jq��sn���|���t}��[����s҄�|U���_�������_Ae��Z��7��DS��VH��'ie{�g�<c�[����~��K�>5�(�L��"888����3!���]:A؀�!���[�@rɠ�נU<ﻌgL7z����Y��܌�JX�����������`Ы������䍦����r���讶jp�s�b�H:�I9RX׼��Ӄ�k�20�x�U���4/���t�rL|j�h��nq�ÜtKj�������6�K�۵��hf�+�,���D!�̎"ND\|<�]�����/g>ߴ�9�6�F�c&�6���m�\��Q�q��Q�YOu��G����^\A���5�c�T
�ߑH4���Vv��U�L@I���3����{��!����N�������_[ز��b����s޹���f���u��i=�l]ڀW��M���z��z�/8B���z��Ȧ��6���JD����r����%�,A�&�.f��w�1�fm@���K&���I�s��m���ռ�#N�v[��4F	�����IT����k(ϐ�s+��C9�^$����ـ��{1zc<oW�	F�M�h?�%�j�
M17lOO�/������佸0�����Uh��`��T1Z���8�:u�)N�I�l�7�~����?�z��&�̓�/,�r5J<���	~�U@���g��9���Ǐl̀�K���[eF��&&Ym�k�c��f�p�s� 	\�#*�i�b��{��K�e��j;%a�:-9/Ŵ�F�R`��vc����('I�)��tɌ�Acw�!3+��	U�Ҫ�0]�\�u�11�� ���(�C�ߘ�d��&q��/Ug���vvJ�4����	��|��?�]���	eӗoBN�~��oH�mԘZ;�WS�J7$4�fa��%C�i܁t<�kJk�_H)o�?ğ���㒂L y�%�Q8��␵�I ���Õˋ�� M)��A��ԣ0�c�^��{p����r��B+��l�0g}Tg2D�ǳ"��մ�Wo2O2|��ܖ�4N� d������c���%E��zΩ��%M�C��6C�Q+�*�pZ8Us�N��e+8,��#�]��SY��s���#�!���ƹ�E ���7�`�S'�n��q�}�
`E Mܯ^׉C����E��[v;��~�Xh�B4ƶ��\���v���qGUY���Z7*�T­}1�o2�k���w>�i�&̳3�T��c7w�+�=��ȅ+�Ȓ�gK���{5L
���_��2bO���K�����z��V�;�N��/�z�e�n���X<�M�t˛����zʠ�H���H�9�%�;xON:����y��Ʀ#f�w��vF���=2^,�.�ZH��C;�Pr�G����[��I����9*(�Â2	ESO',9�uA��t4FB��z�i����2�k������w����H��U���2�	_�r�#~��U۹�Nx���"�C���P�`�*�:b$��諠��>K~M��Q�mm˻�0���R>o�I'��J���k�p1��w��PW��	������,��-/6��;'��ݤL�ryt��L��8�����`8�x��ۃ���K$�ק���׊�/b�PUO%ʱ�_��/C�i��I^�k�S8��/A�Ŏ.p�����Zf���k�Ȳ'�ms^�������J,��'֣�
Cݕ�i?����P�刿*���ޘ�3�Ja?T�z|d����/m�+�k~�u��=�����Ν�#y��x�&!oyv=~r�fU��B)��`i�B0�a����/9�U�nh������l�{����+��~��"��wD������@*_r��B��_�OO�>������%��Ta�p[W:���X��u����u)b���*�hpL����[mlr^X����A~�����fd(��,3%�_�ԣ�����G���P!h�I'���β��aZ@���wչ���g��d5�V�煯� ����3dPB��y"G���� ��C�
�Ę,���N����M���O��f~NȀQ�~~:��	`7�3_�������y����H��u����8+�NxаCI�mE�#����
��o��#�3UV��AU'������+�x\�7~�Gr,~IT��R�o"r�R4trz�m��!^J�.��64��@O�)�2�V�x���g#�wܑ*5���xFhNN��s,��{�_�����G�<o����T��AO�(�vɰf�Q~4��L�h�7��}uq�����tI]�]�-�#�Mu���Ϙ3\�O�	:2}�Q��߂c�_k�j��Cl��|��dtS� Jo�_��n�U�p#+�;�Y��|&���?��b����D�`C=�g�,7�?v��T;A�y�L���-V�Ϩ�u�O�r�[D��>/�;*��AqX�,VP�;��Ao���=pm�b}��~�������RW��ϧ����3����� 9�gY�mk~�m�j�{?భW��T�k�K���h�5�8�Ϲ�{�(�7�7E6'�F�[9�2p�~�c(0�����i���qg���eO��S�h��,@�1��L�(/��B��L�ʹ=�@�Z���h���j�����:Ô���艉K���i�n��	���$��nw���% �V��	��f W��wm�,^-]K��/��;��G���6���S�t�W2i����{W䛰�J&G��
P�{�Y#im�YӠ�t|f&�����q��b�IK�L��BB,M�-�[,{Y~p� �Qn�Dp�4�$$��qp�����жF��
$R���}+��蚷hߪ�w�un�S�O#��M�,D���N���yCިa��V��^���l�����u�����m�F�bP�W���c/�I����n����:!�">l�J9bw�/��������~�k}������^�dJ+��k}1��;� t���"pp����]�¢B�������W�w)�?���h�u��/�/B��d�'`�L��b삵��'����}�x��KG�X�B�nu���W�s��r�*�,S�ZG,X��A���1o��x������&�b�3�ݟz~k�_�JOy�Γ.��5�{%�Q�#�T��C,�@�)�L86eژ^�>t
x����+j�2�1�e���;ݧv�{(,zB���=ݢ�('�G�now���E�6A�����W����XQ7�h\�	��u4L!������0�&̌��S_�L��+�Q����3B�8�p��
E!p�3vz�(�B�9F,7�9,}���i�w#$�=�+�MT*���S.�g.x.����c��ɀ��Ɖ�T�ڕ�BF��e�̺��Z`����ls����R�H?��D�^��R�������� �fC��
~�I�9>�_�xv]�^�!*vځ8�����H���wޮ	����	f�kψ�>�B:�_�B�0��2I�w!X�A�V�Q[&���!k ��P27���r';�E �_���9�t2[�s␊����!��`��ڷ��Ң(}3⢷1��7��x�G�1��R����O��닋{0e7]�Br�z\	��q���﷭<{
�}���K+���������<Gx9�x���/>X�*�������^&N7�q���H�}����ғ�,E�_!��^��0r�p��pl�r��u+ժ���^�dʲ&+�i���ܸ���"(�����o�\�[��@�Ǐ4g��%S�T�#�����Z�Bφa�)lUp�\m���WW�=ƻ8T*��"}=f���}�`[��jp+Q����~�1A��`K��7����0�H{���nw��-âb��*818�z?���<����~�x-�!55uo�,�Y����3>��u��ppI܃��<U���]@�2�?Xc7Dy}�A|I+(�:W�aip��`և�3����#��I��e敻M���N��rï��`n�0����wB�P�@_4�@� �a�G�cv��`I�v
r_��3U_O��B�衈��ɮ5̏�[�Gs!s���m������Ͻ���j��R�ѵ�Ը#D�������}V��\���3a�G�6�}�6�m����F�2H}&�Q�So^T�apdEi^��z��`��|�M9��@ݟ�*�����rz���W٬#ɭnT?��1��'�/`e-�i���ڭ�8�,h;Ӟ���)�Ő���-V�}�G��=�x��o��HI6�x��{^3�.xF*�m�b�بR��d-���n>0��Z4���`H�u^!�'��T���^�S
|���?�eI2�L=�?>��I�;�?�d��i��=�P��##���|1�v}:�g��6F� ¨�P�pj'D�Y�u��	h�X�`Н�S~^��E�R.b��5޹����K؍��Jm	�=�(rs��U&��7�~���Yȴ���t��� ��(<��c:ds9�*�qEL\� �5x�%VF�FJ!q��d���=U��Kx���%�VSΙ�p��[�B�Mk�p*i �$��"r���utD>�.��Ou���ΝKbC B �[�8�Lj#+?V<�Zs�|�թ~f�� �]K�lMiLP���%I�þ��f?ʊ��Օa;��r��a���_�t�,i�δ��+����/շ�w��a%��t}�sNlC���-�
'����� wH��_Ma�nmɊX��^��Y�;�r��ӱ-�������~2N�B wHj>
io�P�*��s��E3���{�g�9x� `��B��:��D���:O�KI �`f�s�;"�R���㐸7�h��Ԥ���40�c��a��9-)�o|�x�ǻ�}�HI�k[v�!�[�IFG�T��M&C���6���Ѝ�'0�w��_-6�}8U+����d-c�:���UW�O�V�98�o���(��b"~�V��K�t�.�C���8��{[���dMV2,�Y6E ��N~�1����7ў��z �G�N������f��DI,$����F�������JO�_������S?v�z�UIbH<�����wa�W]��,W�R_� �U����;K4����=�Ѯ���9oP'FrUn�{�C��?����7c�L�c�:�u3K��i�/����qJ����r���âB#�v˴G{U��b���ҝG��R�Wm���^�ܿ�+,,�Mo?��yZ 1��(mjV�l�.R>����AI�Ej���U��쬺|����E�9�`�b�k�������m�-��r��x����_�<*�U�t�:���$[֬�����]`]��~h��D^��|2����8�C�x���R=��/��/�`�{{���v�@#���^S��)8���Z�[J$��R3��9x������{u)�f��hɦv0N�^����gXH��
~�������
�\�.�^Q�����W?{�1�S���y�sm=IB�;����S��������Ri�N�w���vz��^џ�`W�d��j�Nis��ί��&X�`Qi�`L�vV�m�z|�pɇV%�q���b�M�\�����~q�8ly.�j~ӌ����f���^ޙq���_Q=�D�u�@�<�8ַ9��X��qc�>����u��~!`|B�	�::�/��oħ�o�	0Й��)�Z.#y�h�wA���r���{~�e  0�P���t��m�ާ� .��`��֚diߐg]*���K�����췢�/��t�T�"��h��)q�����RQn�s ��^3�4���zܲ��7a��7��!��9�
�[yڵ),��8O��@2G��~�E��zª��^J/
U��5CGa�tA�f�V�����$7��j�+m��0��wh�~='�*|���Aa��� u��[�l�[ngy��g2�[�,�6���G�C�!�>�B󰌬٢� �DȆkG��Z���=��'��\C\����s�|h�r�^�|�W�A����dV%Ь��)�]���^������z^������837�;"��3_�}��1����/�P�|��#b���TfE=���#N��cҷ�^/�/�h��-�U?P�s6��2�?W/�G�\2��s��(9�VؽU�&��/5krW0A�gy����F�"l(s��"��Wm�v��������W��Mufn9�T�b�e�ݭ�L>((J��+h�'i�ɷ�)����s�D21�6��gRV^0L�P��7���� !�~�/*hJ�C�x�Lab(����7�N�?V'�2*�;R�DM�A������;W�#�I���2�P��#��c#��s\T�i ��5��>��Yת��И�jҕ�0����[�����ָ���v`�Lk|M�]{��u
@�2���p+fE6�_wEdY����\��z'�g�iʉV���Q�hwG�?z���)z��L�%m&�~��6��nz�=�|��A��Wx��\ab����-:�n��eS3�V0��֊���G{����m�Š6�S����փ�v�v����zD�gw�)6w����/�љQ��pa�l?��H�<�|mD~��cj!����e��*h��4i�vk��Txp�&�"�� u�]v�@����$G1|@�_�u}�����c`�X�3�K�� 3�
��0�qQ���l���c�S�g�E�ǻ��6�!�N����>l	)��OkD$��x5o��V�ͺ�<}�=��uƉ�=�ݍ�>�e��]�l��h��q6��uJ���*��yI������F�'�`������0��9\����_H��M��	ﾉ�QJ�u�ؚ���oPu��3OB���U�Mįhu��Q��Z��*`�7ߌh�3`G8M5tM�f�@	gw���Rj����{�0���1���C�#;+�f��i��M;X��=z��cM�P2��7�22}v��x���y>O��������+6�6���b.5�:3WG:R��h>F��:�<o�cBޢ����A��m�lQ����<��Вb�����9C֙c��[ ��]F4�`�}�*g����� �r�6�{�o��`�u��Xe*���N����s`�����ˍ Q)�������{���1�=`v�tM!Z-�.��Hi��Z�@�?��_�Xr�V��Xsň��ca����w�
~�Y���3溇sڣ|1�)*~�6;~_���ر#+?n�f��2HRjs�f�~�`�t���i��Vyc�f�m6g�B<]N�{$`*�`r���h@m0�t�gb4����"2�Z��+u���V�83ժ-`�H�H��B �ZrE&˞h|_m�|�b3q,��I J	�m{J���|9�2{@O>'L�Ǻ�g����$P$���rYf=���7W����Y���*��3�����@ڣ���o�b�����YT�n~�S�vzRC�����dI����D�}� J[tfe#C���mD�-��p;�eXn4J�<�
�Ѹ������|�-g'Af�ӕwj˟�z��|3G����3�v,(��m�#Gh���P֓;�(M����`��A3�&���ai�����W.|M$���b,�J*�O���K�����ٛsu�hw���aA�P�̓@y;�U��W�{�J����Đ�.*�����M呿�HplM�ID��2�f��X�r<8� 8����U�fW�����F�P9�����9��f��ڨ:<DD;���F���y�N]�^`������]�Qk;�P��٪i�ɹnE�}6x���j�*��̊D�;�"���l�"�9U�?۬�vn4m2����cUNڡ�aq��FV&|u|�!�㴓^�Y�j0�."�D�m���������3F���>��~	i�m���W�Zi���!��ݑ��K��|��~��)�����^���U@��f�n��dCP&�'oVT;z�a�`�/:��Q��"n�^�����m������m�ѓ���.���ڬ�H7+���K�WU��Q
�c;xڳ%d�t�[~9zi=7���U^�	�N��Cz
pɢ�7\3d����&����+-��p�����k�_)�pe�ô��y�]��!3k&���2��~NG+��?/�c��x!�8�_�����zedۂ��7t��F�o��Zm��F��|!�I��mqZ�^�߽������_0�%��R�Ae��6L��ys��DlP�e�s��x����W���v'�G��
��%���E����7�<m�����6�J���Z�aw�m�Fr�����;�v�[G�� ��Xެ��|>����z�2���j&�'���U�=m],�~��`uz����VMV	��ڊ�'6g$��,~�x���3u�0�A0�x����M�3!)��sr��L�H�0Y»�Z�x�K�4z���F\���.�A �"7wc��B�#�Xx��7V�B��OҲ�Ϊ���v�p'��63j��S\s���]�ٸ��a&p.6�S�������!Q�]q����ll���`c��J,��'ٶ�
q�9J5d��_��1T]/��ߋ��}I��w��V�;���)�^��Nq���:~hm�G���4�|�z�umܢ�1��a�(Y瑙O��r\V&69�
�	Ӣ2RO�ۮ4�M��ۈ�� :�9�����m�G�DJ����Q8`��F+u-s��?Hc�[�v�ĹF����{����e�@��}b?=PIsP7��&4����DX��:�8�{i����7���b�\`PQ�}H[�qk;j�B��d�$R��[���+K�%a������MfI����&\��wD�.��+zg��.���u�k�{1�.?�1ӽkn�{(Xa��v�f1е�q�ۄ �3�[�����S�'꺆�>dO���������凳&>��Qs�aO��A���P�l��V��O��0��\��<Caa��ᙠ��������`��JJs�G*
�c�2ee�/� ���[����B}��F���"h����R���Vj���J�KDi���_?9��찟O(Y��uTP��)`կ�5��&oV���i�����d�ɰ�_�ʛ�E;�1���e*�^.|�X���Z7�\� �2Apι��x��6�Y	Œ`���\4��fD�b��������h}��˕�h�}�A��B��<V���� ʛ���} �u-M"M~��w_ƌ�t1ߘXŋ5�lF���kDR�ӫ�} �U|����̈hh���9����F-�������ν�/Z�˚����c:�p�e|��F���Y�w�f����O��TP��0W��!��J���=h2<?�7��f������IX�{f� M����lF��ѵ��%�K�m~p>�f��M�$�z�o�J�������-�r,�y>�c�gx��k,кNz�.;%���g/A����P$ ΪSq����1x]��|�J��I�}r ��O� oޯF%��"]u:�P��fƞ��i�E�f��]���fa3?��<庣��wM���z����|9��)	�o�֘����3hy�+�j�TW 8ʮH�Gb�4�U�3ꥄ�m
�,=���j-�E�V�䤑O��!>dJ��&�gI4i��:Qi�_z1`���",��M4�q*@;�9F�Vh�,ӆ6�%Y�M�ɇ�l�{>n5���dp�������u^�7]Ѯ8��ı8%w��J�D(3;����"�Nܚ�f�}��c��1�v[��ؚ�XoL����Ұ|_���5��V�ԆD��uZP0?�+�`�+aN���>V�,�Z��}Po�Q��Y �`ͫ�=3Jm��h����*I�@�����E$^^���r��5|oC�/
w6�����?���[U���(>-د�X�/p���:=�w��إr�:n��ɭ��1��U"y�������O#��H�2o�=}�v��{U�h�1���u�����̵�n���t�����{_ᬫ��c!���9J�f�����*��yPU{���b�po�Ӓ]Q�JT��Q��r�M>�l�D�x{��pTs�4�������A��>�qܧRM� [�9}�X�������$��]1P�$�j��N��u��Z���d~[A���Hk��E��&lȉƋ8�Y��^����o�;j����Жe���&,�=G�G���Ԁ?kϧ����n�ˠ����22F��T�(F��@c���@�ݜ<�/��3*rn��N�L˘�Ծ^�Qt|�Z.Mx�c�n��}�5��?�$����\�e�.���Rd;,iTYA祎��(�vU|������i$�p�	�?�����L)��C����s��\�!�����;����k�qd"Jp6�|��]�4��W~��Օ�|�����;��=��E|l����kU64��]�Z i7Qid�`t�~��|�(6�"֫h�3bڢ��u���23��G+o�<{���m,�b���d �m�j�-��W����>�%��5~�+�Z
#{c]ݨ���JA}#s#�����	q�ɛ΀S��M "�x��;J�*���O@���]�y`����U�*�ӃFА�hG�"&W/�W)L:�W'��G&ï_UR���A����+~�P�h�M�&�1
.������oV�/��Q�-ۡŦYe�%���ى�ƌ�o�$x<(��a^��X{��+|	��L��� ���(;���/_-��g���I'c�%�+�}������נ+`ZO/�}�Z����H�y�Rd�X`�d'"���:�&w��tR��U,�Q$��j냿]3�Y"{M��W`�n�X���?G���2���kߧ<@"���cc�f=4�R�������C�WG5�JJ7�H�t� Hw3jt������a��etר������<���� ���S��������������E����P���x7ͦy$ �kU��,�8fl���P���N��Z:�4�r�$���"�c��'O�p<M�)�]}��^�72u�)����+�y�7��a6�nM��)�������]I ^_閌[k�p����Ki��I5��?�x�ϓX��v"aLr��<,
��������`���#�VJ�}�|0�1�8Q'�kD��zR\@��EK?�Ŗ&��l6���m�Vl��D{f�t]�������+�����m�9�:f�d�����3��W�_�h��H�xMs[���s/���o�p����r�����R������]��]���r9ByjU��|Zf۵�˒  ��+�8 �q8�l���T�]|�t��!��$XH��}��+^�N��lrۇy\�.��@��m�\�k���l���{�*g�����py�8X$^C�Wj1�L��s�	�h:Fg��b��>��m��`���N|GZӾ��������'&($�7u�����z¨��r0jW�8�|�g�1�,4�'�g寤��1���j�c�Q����}jTj��&��e��J�ʎ����^o:�!>TuG�$^m	)�3�C
�Hz_:0C�β��h"* �_w1S��oJ�����
��8�J�µ��8G�l{�'�øx	Y�5�~���e��O������:��>��6y������ː�Z��ó}V���4&|��'�&���ޡ����.����q��Z*���T'����)&��\1	y���T��i�6������ʫ�j�R9xx>�U(U]ҕ�oկ����M���O���F��UKg�U��u3�f)F�Z*5cU�2Ԕo@E\� �"�)�ָ��o���W[�ц鳱JJ�-���Sp�t�f׽%)���5�.EeF��?8��b1дs�c��r�'�6�����\��q�o� ���z`xUO���ه�R��2���.狋���72�}�p�^_�JQr:N]m_��.���习(xux�o�0v�M��+����s�OƵ;�h�jԤ[�x��iȚ����1�� �N��\��̜�P�N)��v,Sm<�9��,2\�/Cs(�DM��nSw������M�n�pH�3/���AMw���(m�r�8�SĊm	����j�5N����&�jy��
6]6n{�}3��~�h�Q��x��h��~�kF6��.�K�v�y:�	�`�Lj���+v�	.ָT-O\����R�#����ݑ/����c��}#a�7,o�ENA1Q��PŜ�ɌF�7�z޴w�z�����@�n��WO8�'�Do��H�g��+���K�3> ^t�DՉ��G�,�t2ΚLQzn��M�J�5[�C�L��%�nQx�s'��$�+;����jmHپF>9���ۨʥuo{�ZG�0���^ݢ�X^���Ó�܇�c:8���
o[�3�'����J���ɱ�sG����3��[0ʩ����_f��8&�wÒ!�{[lF�;OmŇ6Q�ڕ�=�v�n.m|)���l�d�ל�h`�P,44C�H�n�|��w��]�d77��.�f[\�U�W��F���e�~�[J�qfK���ZEl-�Қ��g�!F�PI�Ú�.색.�˦�FUZO(�hm�����t�(���M���%:
dQ�㨝�OWX�>M1���A�1�Lul�����XF:Cw��i��Z���<-o��gy�x��c���qe�A��?1?R9�������y��]j}����.���RXi�����/f��h�|���VB3Qo����������|�������h�I��,qf�Z+k)��7�T�=���f��q�\�1�(@t������.��it9��3�*멼��J�x�B�?�������^�<)��/q�o#󲻀����Q+a�)?R�DdZ����'�T�B��D�C�bHI�F����5�M�4p�{�&�ro(}{�ǁ#Qs��-�Π��S�������n������� g�r���$�>��XJ�L�ߢ��_��
�����^�|?ȸ������f~������Քב�Z�)�G�Hqu*��6FR�R�	�{�R��dL��a�-�V�^�R�X������93���US)ͤ���횄U		����G���cVR®��]�Vwvl'�R`>�o�pa�o���[�kT�3k�6��8.�m�?>%g�=cKEQ��\9� ��))x�$B�r7a��83;��F:'���r��CY��J�����WR���͐�c�FYc{������E�H��c�P�T��87@����-%�y(}��\k9>��\_=p�^�g��!G��S	��x��w!��tq�����jK2KwnR�>���tz!�*��8��b!l=^�l`O����K\�T�AN*��pkm,�����
^EE�	����n?PTS!��vO��lq7�����L��_y^m)�a~�/a�:��A��;_���{��=�@]�ۻ��Q%���w�G
��+���Ej̾G��ݭ^��5=,}vH�L$뽔�D은��[Wr��/q�!{���	�`��yː$�y�M,�M��Z���	���@<��5�t�j�}��H$ �`>ʁ�es���#���?���;�1�R]6ko�#������
��L�'�M��RȒ��$ZW@�ߙ�T���J�Nc����!4�<g�1�l�<�>�)��M%�V0�SsedZ��适�l�݋�V��`���u�ci�$l�L�5K�gf���i��.��
��5�� X�!wG�����Яl55\+ѕ]�C��$'ְ�����T��JI����:�W�-��4�\�K5[P�{�\�)�)�*u�tL�BrD®��h�e�j|����*��~�ߙIP��iH�]B�6�$F[���#�&��pi�T.2"/��h��5���?y��T��o�Z��z?+����*�&�PB;(J����#m�&��c�z�����7>\fS�����F��TJ�~Ytr'�F���s����Ϧ�EoD��Kd+�bh�t��<���L~$���YU��^1�&D�xπ�K�c���a�Zw�9��w���uA�M������?�-��騮��U��&S��WH��i]֌կ���yW����G��=�1Ò����j��:���P$�*��.�� �_������aZʤ2l���|�}���?�oV��~猝S�tP�����I,�UN���̼kM�O�S�-;4�(C�o+��_�{1���(��u�I�ku:�i���t�P1b���)�sI9����)��b��a5��V�/;�.�w2ͣ.1�)��Om���c���4��p��D���xG��(��Fp����e;�v"�芮ߙ��k��V�zQ�1�9�8pTT֜�����/���KIج*>��ƕvHkp�d��d?T���J%�h)�%����ˊ��<$��΍+��Y�t���Qę�]��g�g^d�a�h�L�0ܑ���\<��v�0�_�=�bQ9�K��N�6v�y��'mտ�tSV⻷�q��Ч��cG+�:6�\g^�44�#-C1��;5g:��&<}j)���]���I�r���J�]70x�pu�����`"k�Iw(gv1�ss)��3a
���t��4-�X�Ei����:IfHcb���R8��ah���kTʆV��/}�B�#�jLdQ�!�����+Ȉ��7͑�4)��U����f���T�)�%ٜFY�uh.�o�(��]�g�]�nƻ�\��!��fe�$�7V��A��q�#d����Q��ȜZ�a��o�L.K���b�V��J�:q����h�/).����hbC���t�MZbeOE޺�mm��7�͚W��c�W�������o惡�3}�_~�oi�K
���j9���L�8?<���9%}�mr�(�������;���s(���$�`'�ojzJ��BV/�<�`��cy���)M���Ӓ�;�5>��HR�uD��QQ�L�is!~����_h�m�*,,���W8��K�86�zc�� ��O)$$4��lX����	r:����������]���7)��c�E���?�_Dn#*�Xd�X;���}8:�f��_���Ӆ��hE�q:V�i��o��~5M,咒����"�!Q�9s��w����	���79suWo5� ʿ����nm�<����'����LE�=���\�ߎһ��(��~����1�z�CV�׃7�:�!���ͦ��� ��d"}��)_A��=���i��V:ڧ�mĐ$*u�ۥ��b�f�3�`�W���6�uΔ�c�iQ��+v���$�� gJ����:�� K[z��Ո����ow���|{���Q�x8,_��"#�V���,-E]^��yx O�{u��I8~��`�T)�g�������]��)�+J��\�LE������ME�J�(������Y�B:��K�?E���N��܈���0��m�.�.%n"� U��m:��r��Y�zE+ZXR�b� {ȿ.��2yL_b��Wۜh��Dc-� ���,��Á�}��ޒY�N}�|쭰��H1�,8e�l]��|0ɌeK2m2�'d �
�^��[j;�N0��|�њ����<q�Ӵ�ץ<�c���a��Y�s%��MA㇇22��Ǉ��LB�¬��Ġ��p���U����O�c{8�?fm�o��߭���@��v���v���c�D��65�����Ԛ����[T0Hs�r�v�s����h��-��A]�)xgB�Ӝ߇A�Ҡ��B����������/�7A�VP�Q<�ˌނL�&�֛�6��@�CTCL�P�?��'���B����ǻ�X�?�R7YΌ���J�u�������������CF.���X�eXF�;G�#��T�b�~51oN2	�J~X�+�G4��]5���?D�vD�1I�I�+6r�v��|��^�TԘ�'����p�Όx��=B:1��P�_k���/��V��h[�X����4"?��Û�e����x4�o#��<ӈ�׻VzJ�>��;�qQ	�c[�f��F-�'CMv'
tZ\��u��j�Gj��c����)�ޯSb��!B\�{{�/s�O��ͯo��ٚ����=�&�.�<ZN��{��De�yOO�u&ɮ�K��<�r��^��:��±�������K΃�3:q��q��FU��o"��x��ǭ,�s�V�@WN��0c��w��kJ�b��b�P�$�I��7͏���M�^]s��{;���*�1�k�|5/�wO�_*I���&V�G}����3�Į�ofW����#S��+,��H���R<�=�����L��*ɭY��y�n���q,$�Ǵ�m��Qq��eb��z�|bb1���;��H(׏���F4�3���XH���~G�;g��-xľg(��'ԙ��E����u��(�ɏ�D�*am�~eM�< ���fa|���^S�)��*S�ovG5M#zB'���K��'<�����uk��[�L/�i�(��o�����P%�������t@�o��~���O�km�s,*w�se	u��qܦ�9�ݐJ�L����fMs�v��s'�� �����9���e!�PIj/ن-�Y���+�1a���dok'�.ҫn����v�������y�+d�o� 	][[[fdb�3<�hw�K�zħ�Q������<5�|_f�'f���heo�����*_�0]����k�֓�;�@B��/�����GW�>��'�=�b5)C���3��7��5O��88� 5�s�g��Y�z'��Bx9LY32]yق�@80�m��#�|fE�Z����.�YP",���$�u��b���)�gS��ͩ��փ?V��j���&��xȹ�ww�f��/x���;���3��S>��U�=*�L�}�j��f��=T.p�{vԄ:�}�]��)���$Z���yc"���JV��ӻ�H���1yL���G����+.a�K;�Z���� bCm�����ܺ�:Oں���j%�3�:���kFOFp���ݙֲa>h:|�~W0R��ıe�+��bg�?���+yi�����]f�ڝ4	��c��g��#�g�������W��N�AgQdJ�k�<�1�D�E?�:%e�9�:'O��_n�%KU�����ͣ�K����r���+��³nw[���ĝ(���3��p0�뢨��iݓn�'�i�R�k���J�%�����==�m�ݲ���ݤm�� ���z��G[��������>Q�=zYĭn�X�&]�--�-u���#z�o��|'#���n�Q���O��+��D���n�޶��5oaW�EȬ ��ܵϓ����.�����"�gS���Yi��^��6U�^y�b��E�։05n�j�..r!�BBV����X��=ms�S_�q�*�Ȋ�#�q0V�Df�G�*??��i蹆�!��x�28svNb<�`$5���<�_�C�rV���\Z����e���+f	*؁����f�59l�0� Ď�{��p�I�M�fo���{8�L��O������d�yZ���us۾��>BԨ[	/w�@��R�qI۔ lab�ͷ�n]������Xs[:��H��8��h�z�]�k��L��k3��&s#Zs�I��i�"L���IO�d��UP�v� Y�䀄� �˹������ϱ�,t���r�ړSU�'***���s1?��z.��d.��u6����	�e��6z F�X�L����:��.,N��,Q2J� % ��]������K������6��\T�PO2J �a4kb�*ۚ5��2凼��5�á�e���>f��ݢ��|Q��QNe�J���7$a���ݾU��>=�]ԩH�y����D��7�q�/e;�a��۱j�	�bd�ܛ-������o�o�����N�;)��>��N9�����!�X�K�ղ�k�w�^��z.M;����,dIl�^9]�g�"����?���Ug�fY���7Bp�R1�1�}}����1�ʃM>PxrT�S#Zg�\���1�ǲ�e�$#I���2|Zۨף�p��R�P�����b�^�x$`�x��7k��}B�6����U��>����Vf�񎩆II�i
J���d+��-D��X�>��j�r:?3Qf�WE�o����4�2R���r�M�z�%��kl���tT�Ln��@���c7�֠�C�E��--�X]u�im`呶RfQ��H�ӯ^F�. �e�-K�K	5�)i-ؘbbos���e������}�j\5	)ά3 ���2�%��X��(�e�L�����6N��5�v ;��n~��Ԟ�:g����]�s��bQ�z!�jek+���M-��I2Z���|8G����fsd��k׳�Z���3�'V�J6�B��ڿe[�Y��G��$�<�����J���~T����qs)������\`E�E���;���@7S���x�5Ԭj�z@��?&S3�,1��z//u��5��b29���)� ,��m(k4>�-W��?����@� �B�Q� �� �9k���k)�� xIDs���+�Bd�j��^�1�0��WL�#���ⵇ7L����`*eІ����$B�q���DnO<,0�������>1��ӣG@pۨ�k���ͨ�*�Ͼ��pQ�Ȉ�C6��==�����!~<�G!��/�W�]�ɘ$7��SZF�j�H�r��
Yy��x�*.�7\q_��|"��lC���-wd�,I�]K�P[��*�Z�C��@�����e����O��V湊H՞_ߞ���9BA�T��o7f�	G�0�X�b�)�WCufM�`.f����M�:+f$[6|V����ԖAf=go9���?�{*N7��me-��$L�Y�C��!�?�Lt��'��hή�Q�
t�o������vՑ���!F���L��ηY;���~�yUU2�(�QG�����.q�%�uq\�[]���:�t���?�c�k�zjv6��MtMF�
�?ɜF}��h_��擐<�����������$��JJ�j�^�m}��J�2ś;"�n~�`Y����>�l���Ǡ�WVE���iԅ�]2��pj�\}9��^n���Ӑ�������J7���z�=N���j�z}Ǳk�ʿD�ӌ�G%:���U�En�uq�������4���
����qΊ��3k
�:�w�Rm���#���7�M����i ���PV�~n���́\I')�tuɼQ
~u�UQrn�~�aP�RE=�h׀��O�kG��r�yG:'h199)�s�vy�L6�~EHH�st$͑	���\s��:�9'#��̴崭/��GQG�aW�>��/sS�4�Eϋi�ӫ��+�F;�,�-�E4(?Po9z���;����k��U�Q�&��K� �����7�⿿[O4A?{�cy�����LJ��h��נ�&���4`'�X�y�l����?v��m����K����::w����1v1ȿ�KSuc�^sN:Q`t�^����hp�g�;U��*� �^΂QJ^�P���l�C�G6�ᵳf�T���VqAW�EE�QǨ�B����Z}�9���������QQ�'k�sm>�#��a���<��� -S: ���ηG�r(K��i9�fǕvj�Y4��
c୧Zf�9�ݟM��e���S>�[���"��� �Y���e&����d��0���u��݌g��R�QY��r��Fx
ʦ���g�MKELP݉?�z�
�$��M�l� �RK$�0^�/�LDK�� @����~kc��j]�}�b��r��&�0�+���-o>%�9��{��#����]��L��{qw���A�P��C�yܧ��{�t��0ʉx����D[�0�_f(C���|Qp�v����۝�\!u�>1����++c=�%�������WB(2��HS<�U?�vEEE�\��K>����u�yԲO~Xh���֟�������a�2���,�b������+R'A��8ݹT�۷���`\QXN�rR�l��): ��|0#�>`hͽT���:��p�g����ȕ"|��_�{2����u~��
%	
�!����u���VF�Z��� 
iTӞѬ$=]r?j� ��F���=��b��w&-K�T;YXQM��z�,�]���?�2�b�`�e�Ȼ�`>�Z,!��mA{w:ppp�6���r%����+++�F|B�,-��1K��У+����n� ���+ޤgd�� �U~8EJ����:;?��[V��s���_�s�g���_�W��K��T���h�a��T�)z�7*a��K�+�ፒ��T.��%�)ed�h�2Ś*N��/~_�B��Ő{)+p���G�>&��_y���s�-���$1����	�N?�a���
g���3�w�9X���r�����RLy-�3�2���%Bs=�+ѝ����8���B@�~��.�D�m"����S/'Y��Je�|6����`�jV����/�N��)Y_��B�VV/�Z�0�.4�f�'�9�WJ�nR�|�;���IqHm��td@}^��Ld��c�	��t\�7�%x^pWPT�(��N���N������%���Ъ�e�梄xA�ǟ����DT���Y�.��n���trp[�����R.ϯ	^g���"���-����5w��-ETUN�$BmG5�W%O���3�!g�����	l�Q@�
j}�{��o��D��_4Ĭ �Y��V�2��L����/[If��q +�����n�޳]�T���n�\B���m�vG}ӡ���OV�'�fB�F�2{�~�sڥc�k�{f�Î�e�� QC�O�*3<��ڜ/�>#�C�p(a�ax�uu�������rs[M�7�`@H���T��#T��e��rCEѱ�p�[���3%����5~�]B�d�ޘ˟�W�|/'20���
�Q$���	#9���p�掠��\o�H��&�N�9rAH���hIZ\�W�u:� �ѱo-Aϥ�Y?e�g��b��.��������zk�[v����R��7d�u	�n��\:US�A^�����&�����7קb���)�X��nA�adF$'mD�� .������F�֪r���f�p�,@LU���*j�ev����50ŗ��5�����<0j�x�ǎ�aǓ�㜢"&bӆ�����p���S#$�����_�Y�:�Iu�v�q�傭s�Z�E�Ď�*����I��vc�iPS`M�fH��`���DV�_��~ǡ���;i��jK�>�M��{���
*��Q��-�x�ڨz��W���J�?3�|Ye�"g�$����+2{hll�Uo���A-�e*���4������oh�oH9Fs.�b�R�n�I�.j��֑����K4�4��K�T�d��(��e��T'�^n��7�3LY.wbF���z$����B֚�ۣ�|�p�W�B���rn�l�YhI=����w��%�!�{x�xy��b��'HW�#0+9�z!�7��U��ǫ�ظ��fh�W��h7x�F)��lӲ���p}φ���[gm��d�0B��P��dƢL�[_;�l�'����J�P��g�WĀ9S'�N-�?����]�m^�%��6� 2�nQ��n x(j�+�qln�$����\v���Luw�,m��P�L��� ��"�f�h�4Ɩܵ��7b=ݢ�)O�^�t������R:�ǣG)+�۠�u��<���h�]*:���<aé�Y
���$/{"����[,�=��6����|,R�#f�>-2VnQjh�����>^�c�kj��x��|���8n�N�K�z��FQ)H�Pr>�,7��Dwt�[|B���̄�M�e�i`���P
U�,P���q3v�+�&� @.�Xr����0��V�'��4w�a�BG�4-�^Y�X����9"�G���~��}I�V�̑ +��P��@]�9]��&�	��F�'��	##���V�?\�X���yE�������\�}ʨ�V/찊��T��_y&���]��/�1_X>BG�+qh�	�L��4��O�1��1��b�X�P3�n^��!�E�=�����_���l��G��6��Lpn�su��=*����,_����O�yU�Y�4�ߣ謴�̦T*�@9�֗��B�&�g�"�>��I<o�ӑ_�2~jF�ڿ�m7ͬ��}��WX��k�ƟU�ig��9mB��������(�v*�PX�pw3���^>�'�?6Q|
�{O�g�%�H,?�H���y拔	� 2ܿ['��H��6�D	�d�^�ip1옒�Q���X��U�
k���#P�O�+��u��:�F^�n������z���9wQJ�+�G�<b ������o'vy�8��� ɹ'|z|p��?�7��n�B��~����Q������Os���={������G�V��w;qc��û��c�>�� ��5�U䱇;=�Y��9�p�G.64o�@8����e�V�%ͤ�w�S*�o�����
�~�d�i$g���q�3P�����c����I�$�3Q�Ҳ�]>O�HF���3�:z�h2�16yT���b��Q0Ks`�4�^��6��N<�vʞ�0�I�QFY������OA��fj;�Fa���*	�k���)g}a���wH�C�j1)5j�f��EE���z�G�`:y�R=���� ��u��h�D��:�/�K����n2�o�
�N����1��vP�zSX �C�e�Y�~�'�WV��?m�sҩ�lj�Ɩ�w	
r /�?��@]�H�1	��6N��+XM�z�MbiKyU6���,�s_w�,����7��\6�R�4�{Ґc;b��pµ�uWo_�ؕv��P$f6�wm�q֡Ƕ#�(���k4�.`E�jW���.�+�o�&̔�m@�6}M�(�q�n�uM%�r�%�s��˥�4_o�RKh������2�~9�Y?�wl���ʚ�\���:D��O�Pà=.-T�4"d��B_4s�#�F=/����Xԩ|������}6/ظ�} �^=x/ٵ������gƯ�>;�_.d�|�-&��p�;�U9�#���/ID�mXX��9�MUq\,NJ�%U=�(+,�`�PBR-�	����R�����J,}��ޟ	��A��p����݌])&���sE�'�$��'ۊX��	�nOk����Tɱm*�C��@��|��ހő�XK�j_j��8W裆���1�:��������	2FF{!��ح��E,�'Y��9K�;[WxL�0r���<G�a�����2UuuB�p�f�*ż�j	����~w��2y�����i/�i���_Rc�S��壘��*�&��fđM���Ԛ*�DF���h��%`_̦*�?L��<G�	���p%cvԝ��i�b]�qU%ݩ�oK���Ꮨ�y�ЛF��J%O$�ɟ���c��R|���I�>��I�^7�d#�r��0�8_ ]W���zqMz��+#?d
~��4v��]ֻ��#)�o����2���T�P����'����} �;�|����2��=�0�<��'��U�֟R�V&ؑ!u���ʘ+�Va�}��y;��$ET���e�u�ܫ���@)���"�*S��ts0Q�/SaMI	�=\����N�υZ��V�u��fl>&���7����1���JP��u#�?��xP�Y>��G�i"e����%�Ĺ�(l_s�ۼ	�������$�L}��-[X�¡�������c�V�@�6bP�Y�L����nꆔ�1�f���׮އ��k�C+�;��<:�^����r}��U�0^:F���B��ݘb��(<�qj{R��ǟ�U����YiKU���Z�r�̎��8GA��Hˑ��?�0�����oBɁ/���b������z=�����|��#V���/�w���9��ǋ*�J��s2�݈��y�}ք��..=��ܗn�V�fC�P�;��Ne���4���3^`9/xc��T��@u������Bd�L�	��_��oњ��O�c��K��j}r��j��wGӛ����k�N�����.B���*5	��Z��;��-�0���n��(1|��\��sަ��e�-N�hP�[��Բ����;�����r�,�x�+�-��d�Y��剛��Pa���B0��U��o��*ඖǳ*��j.WX]�L���׀��A�a��S�8]�=v�}��2�g���M��T	��KȤ�� ����#��CW�v��js��.���������s/����� D+ς�|^o�B���/,���J��kUO�U\������:O�U�+�HH�1�f�^&�s�t�����sJ��.���J��P��D��oTR�c}�0s���ڷY�E<�J�t�_u��(��/��2�M+�,w*�*��c���<��K��������L��I[<�s���Ĕ��:�Oa�e�"����3v�F��Qx)�W^�5.��<;~)�Q^Y-_C>.LhT����6���?T�rҨ����!��S�&mʸ墟��+��z��Yv����Ϧ*$#���p!1���Zg�x�m�-i����|��ߑk�x��R���b����q��M#$��_�X��qJ=�����`��s����t���ÿI��L�u��9�-��_�[
xz�k�%�����,�+��������!t�vp��A���nX��ʑ�i�(�0u���ٖ�GDuA~~�%*$�U��:�F�%�&�$�}X都n(�Z�Ns��Y6�x���5"bf0���*'YD?�s��q`�rR�؊��]�MQ�rP��
�+�bl��*�, �ku�yI(����)�1�w�:�7!% ̿8&���iŒ��˲�JM���KUc�V}>~�o��1���.�3�����6��Q�FX�/�1�K8a�����yqL�xh=�'͔�(1�k���l ��qBU� ���o��xxx,m	B-�
��Yn�%�f<ll��կL�5u���O��\d�vP��͛I�NOWpT�k�$v�Pģ̤���E'���s�Zx�Y2.i�q==�z*:n��LI28}�M�N�n�at��eiϧ|����ݙ#{V���l��ˋAߒ�_���Q��!�e��:B�z4���Uyk�{n�m\�{Ӓ��6r{k]z�b��p���ݟoCA?K�"�g���0�9o5�z��Ёi�����_�E�eU�'�i�Y�����ѕ�U��`*�Ku��2� �r���R���� ��3G.B�� �h�VA�$Kr����9}�~T�@@��e3�?O�t���. C@�� #S��؆����>�HFm_���r%!!a�\*�\��9�p�ך;'(:h�Z�&��b���p��3�EW�7��������[F.q#a�}��
��#��d��hH���xrM����Ee�-f_��+$��l	b�����[�Gk�߱ؾ�2�����Q���T/A�au��ۜ�->��A1��q�P�r��~Y��g�Bw�ׇRٽ�.�,���P��D88"����s�4����%��b�ȑ[R>�!_�ˍ$5�K7;�'D�oo�p�$n}�&	��ɒ^d���_��jRgP{3�`5���>W��4
���]x��zOQXt8��J�*��
p�m0���j$��('�"�	K�p�Rs*�ɧ��OsX�$-_e�N.E�>�d���������z^����iI�	�ec�oĮ�x�^*xǨ���$a�#�x����E�L6�ȋ>��Nw�M������G�`�r���Z_��y���[^�J׶d����a-l�l�|~�QZ�o�PrY��7��y�-�΄���pH]9�;hI�v_�3����%�s�H^A�{2J=;�?<�X�Z�;[jes����g����vgBEXӒ-�O?mw��0�>�nH�^ck�G).��V3��A�?��a/^+o�:Ln⻨܎ܿ��ދ����� �qƌ42>&�t&X�G���t|� M���ء�$�
?kB�-0'Ek�&0^;��K��ca3�8ڰj����=�Vy[���02Y
wY�k ��Z��I�{iaq���a.ka�-G2P&�yU8�[���V����r44�Ν}���=M������)c�q}#�~G��zn�����.�O��r4�wRY<�L��1��3UF�a4�/=��1����l�������3�f1�xu�	9:rf/@�1I��3c|�;��٧��T}��o��@J_�_q��7���F�g-n51AE�b�Pt
v�$�uҤ*_KG���G/�"����ZK��c�* oӗ�r�����`>f��b5\S�R�E�خ,�� NҚӚ��-�=�mZ����pm .��	�+t�� �r�7�+��aVbv���)S�)�y�Q�9�����E0dZ$���jQ>�E.�&O[�pD7D��X[��:*��A�k(.RH0ː]��� ����ؔW�4ZF��[ovth9�p�C�F�}�ۮ����ߍ��p�,6Ui�"j��	�[���Lϧ��F;� �3�8�����`Z'�� (꺇I�[4%���L[D���<PE�I�:�\�Vtm��"��5Nћ�����P�1y-I�d&��b��
�k\ͱ��Q�<�Ys�5"�PŖ�g�3�-;Kܣ�N�qZ~�I��,_RIObv[�9��E���l���@i[@_,�^ٯ-V�����t.��)�@�Q
BӁ=zW���g��*7Q6�<
}�M�@)P-��᥈3˂pQ�y�ݚ�=A���	�rw�)ǹm�,���\W#�\�����#�1�,����T!=��-#G������}��R�?�w�W��5;��;�7�	E� �,���%P���u���7~gOO��0j�*���H�4��M$!�dh�^,69�  ���T��x������n|����㓐~�&����+t޷�>wp�ȏ��}h���5),e[O����_�[�n�C>	��Zvx�f��tNT��t4g����H���� o�Y�T톗��׋�IL�ͨ��T�]u��\㍮X��S��R}�Ϥm0�J+��p���m��SK�C!3l�i&�KJ�`��MĶZ����E�{^k=�~��B'T�ƴDQX�Q�M�+�sxP�����{���s�y�m�Wk�YMt��v���T���Ȕ�#�(�f����i���>�n�a[Ĭ�%���Xv,$���_'����0c�`���]��/z��O����yw��Q�s�/$,|zҍ��}��B LR'�:5�rϓ��',6ւ00��g� �H���s7�̈��קq}����86���ߕ�t��>F4u�.�('��y��Q�?_�(�[�P�F},��ƹ�+o8x@@�\V$7���Tn� �)}�|��?Ѵ4S�ĸ�����x6��)�շ�n۔���R�I(o��*j���H?����<]_V��;�PV̅0�Dq-N����.�fWԐۘ�gq��N�U<��	�|�$϶��9�p[����hZ|��J]n`0q+��+���\;���X���lPUvww8�"�����T}�C�q�-
"J�H���tw*�twww7R�
�҈tw.�RK/],�4,�����{����<g�93?1�wDy%�sB�!���_N���0:��3�E7��#7��<�\tDD|�LW������϶��K[((,zMA�t�o�
m��/�Ys}!!(\F��:�c�I|����f��q,@aW�x̜�@k��@HZQz?佛��#Ƅ)s��77RT7|�;�K�R�!Ѝ��D;�=�h�Ӏ���S{�U���+�8�^Ҟ6������s�w�D9y{A�
nfLA�����V�a�>��w)���'��֊�U�oO��4���/5Gĭ�g~ZK�V~W!R�l��{y:kU��*`vvϒj̈́��Ī���S*��-./��,
�yR�Ӊ�M,ʥ�ݿΏݮ��v(�a�*T�f�,�/�GkZE����#������9�r~��*z63~������*�jK[�����"p(��L70�wZ>>��yDz�J��X�i���H�W�f1���?�6��G[PM�NG0$�sV;��|w)3{��n��~�M9Ż�j�@�y+)����}�]`cW[����)�'��$6����is2�J	M�G@Oz z�Rߝ��+sC���B����%���Ϩ�5j��)�|fZ��nhxQ�R��k��_��'5��XC<���xt�~�/1���╯]�h�4��v|(m�m���5s$�g�yL�[ηQ�r
Oq���O��?=��T�1�[$���n��6��'8���c�7l�PSS{�_���϶�
|�<nέɅ}�^�Z�Ck:c~����ȗܼ<� zՅ{<)�ڧ/5AJJz|H�쮩��V�r8^Ǵ�-X��3�ˁ;�G�M�eБ��S���z4���qO�ٔ�������ķ@<�	`�ϓ;�,_ ��F6k�H[Q�Dh�c��+M�K��i��ld��rdn
��8��)?%� =v��)>��*�σRoڡ��i���85}G����W�1��Y������qK�E����tfZG�h}=Vn/\���f���D3�S���5�Z�n�B��(�̱��r���^Eƍp?K�������ty�+��k��RXb���"ؾ�O����~~~�l���J�6U¾�kҢ7�K��++q��6骍��5�����Yz�u;����z�G_��J��}̌>��!V.P���;O�>�4��"U�����Z����`�Rs�;��_u�ou����Q�6���r=�ij�=���/JD&�,7{�c�8r��z6����ɫ7�q6��4�E��g`���\z��v��ٷ�֪�RO��x~�Nza��,g7j�qhM�k�ժ�e�X�8�K�A{v������{�m��츑�����o'�#<���ɶs�ڝ����8���h�z�s8�LQ	W�f�����H;��Ǵz�d�W3jV��F̵zsN�}7GԬ�ZKEzd��;?�8|��}������M��y;"www�d?��!�lw��?ҩ͞S����h��Qv���V�i�''�CH\'��?PV�.:��������~�G˧I���|���k�ki���c<��.�
Zd^q��UO$�i�	�hX�����	n�:��V]B9�SM�ڊI#��oz��+��~ש,6ֱO*��Sѥ��͘�llwEK�e�����]c[�$���.���nX[���D\����_t]��{N��?�.	�SV�-�@���W|[�8�1L��#��؊gZ�\��ݿ�z�'%��&!!!|��X<��m���9R�β����i�Y�����������`uu5"���tY>{�eZ��U~Y��)s%6_T����Ö��Q���H�]2�(�@�K޲��+��c�z�
�ml��3�n��W?�QW>μro��`MRm�%�����G%��l�7Kb+G�kN��z�e@å�'5������d.����}���]5��
4���Ok;]ў�dpf�X�[��,-x��\U�� �y$e'�O�3����r��q�w�s<;�uxǻgB9�ά���[���6O(9���ӵ���^�2a�3z����P��m8�[B�2{1f�u�<�Ս��p�3u_3������<��w��J�iii�c�P�>|}�CL�n��=���xO�?<G��B�0uoS����t!�R���\4��z��ޓ�zW?�"�
9:�-���x���U�V��g�{� ��H��� �8���֢I�p�Ors_���38�Qܵ�a���e�$��aG�L�i��L�M��R��i��ڈA���ଂ0t�j^c�+�=��3�ύ�S�����K'��so�frF�zg#�;w,d��v���;B.����6qymf�|l�{�Y/�i���ؚ�JŮ��B������,���Y��r��vX�!��gG��Aݎ?���o{z�F'3Dl]�뎨+*/���ʕ�\��r�w�蔧8�"��+S������/K�_"E4�w�%c��i��͔:�b�&j̶���*c���,�Km$����!�����G��dAr:��E@L�$/tH��b컆�b�`GM ��f�g�͍닺t���3��H�r��$���k��vC�`7(|Z���#��jF5{0p>��~��_�E����Ѵ��lp㮷f�vy��Ukn�0�yư���ݑr=�>�
�m��S�);*ß)���ߛr�K�B]-���Ғ��lTQ�;	^)�%��>���oy��8I�K
��.r~^�0F�S�O0ز�3�^�z EE�cnN�_;���.�8��ߍy*�,��D��
6�[|�\>�|�����g�tu�J�SQ���>GD��r��yd��`����>����6h^���p�����x�>tt�� �y�R�ʙ��u�R� ���$��M��\y�a#��Ǭ����3yն�d"-����(uJ�d�]��R�g��1����L䘎�u����y��an#u&e+��s�''���?��goO~��=�>X8����σƼ����y�\�j�"0�XA6��R�DO�ܢ [2+�BQeO6G8��sa�R�aO<(-�_�ԧ,��x!�S�ozMO' �]]A9������l{3�>���Go������cV1�mE|n��7�3���N�D���B�߉�OV�i��H���v����ӯ� ������G��?�1&ES�>��>b�����ڣ-���UUU�g�6Q�l�W����3��?�0J;�r5PK�5hJh
z��u,�~���a�t�nX���"+xdN���\N��M�,���ٚP�}����Bo�8�\�4��W��7U>�72I��?HڜwpҮ}Wrn����P� ���F�B�5�r����7�\�M����4x+eæ��-��e���,mg�+�/�Jй��N���wL�O�ƿ��5~�5��3F(��AJ.�Y�b��N��!�U�PbKn'����G�āh�^�� �9���ʦKs�p�� "�cY�d�;��A��閱�}zJJ'���F�ݏ��TGW�dW1�433�7^�R &A�������{�]��W�	W� �￈ɪJ�kN؟���b/<��X�&~e6V��6���,ث3��RHGJ�������߲{���Mz����QF�I+CcѧmU+���i�*���/f@�=2�a��l�v~�&��x�|��L�6����wHF�6ų�3���g���$Յ����7��b�/�4��o�ҧU폅c����`�y�]����Kz�/�Ths>j��B,`.�Q����w>Y����.��F�`%���H�<G�g�>�Mp���_�G�e�:���B
m��躍̷�O�l[O�2����k��t�@#��+C����/��d��j���T�"��`m.��@��/�������%�K�S�k�P�F�0b}X����d�E��[4����ŀ-�~�<�6?�?��(�b��O��GT�Z0���K�T�껀 se��]����m�ve���l��hh#{ 5b��:j	�i���)�o���؋�|�#W�n/�R���1{˧��|�m�����c�����Y�X���L��8�?�5b��s_==¿y�yd��h:|*u�1��bǊ;�w-X�Ǻ�R'qS4��!�B��Y6vC$J�ƲE��hC5z�e$�+���ES�����~�Z����U;�?��
�Qԭ2z�p�H���^��[��ڸ�5j1W5�6��2�E�9��~�Ǭ1�[��O@�͚7������01K�
&1 FR��)�ȹGDǐb>t|�Fƭ��c� $挠4
���S��3�"�Uۇ-Q6^35ӗ���ľq'�c��f��墾���D��P,4����-U@�S��T)�u-�KG;�N�p'��(�|�k%���H�	(���xHG�����(9���a4`�tF势~��v���w�k��/�20J����sYw�ah�g3�?���?�p���d��?����tl�0�ő��]�������E�i�Κ 9C)�̨��f��6���tMĤ�迧ZT^K#
���K^��YSjI�0Q���k`�Q�ŝ�N^i&��ޯ'Vσ�1�N�.'��ݎ��tE����z�bK�)~�s��ք�8�*aX��kh�[LzH�ſ�h܇���`�ݼ1s��<��v$�H�t̾���[���ӝ���1ڸnq�MYi������,d�=�-)sUw�R�:�n�$�_��9�[7sZ�^���9�j�䡢8�������U ��%�UXed�z���hɅyE�z���Gq�f|1i��-��2�?5�9�8'^����7
��{�Yg��$������ʻ3�N��cg���rᵟ"�Cq��q�����D�6�u}{���
�˶#\�H15CA��Ws`|�z�O��9�Y2
�z�b�����&�6�������~P(T���o���ju%^��&g�F�P!��I��l'��at�O.vd��|$bXp�ƶ
#-m�H���0�Om�؞ .�,=[���$���q/�(zZޔt��|l�]	�a�g3jSI����.��!���Bc��BCN�"�y><���b�K*�ٜa�
�j��JDM���e����a�V�c����BJa{�&�p2�z�(���VIe�SI߬|+�AE6dF�a���6�E��b���v3ٜ�c[�t����FIOOϔuG��M�~J�/XZ��(|�6�s��ѓ�0�*�|^�i�/�������4�u�V �z��O$g�!ʳ��߶�f��׶ŻI��1�u� P��&����]#R� 7$2%�$�?U�vy�����U+�L��xG�ۧ|���GZ'"@��A�f���� �0��&���NgAo��]j�?�HL�PՇ�L2�pQ�S;��Ɣ@h��C��gP���=��C�
;h�5w�f_mn#"t�|�)>��b�%܍��y`H*������U�!�ֈg����n���@��i��;��!ތ��}с��"�	��h"V���d�h௨j���x�G��+��q8�����Fh��NjA��m����B'�_�R����Fs6!ʯ���%HY�D�Uwz����� ���z.�D��0
-g�cy;<C���Z0<�ŀ��ş�g�"��R�M�.X.�ü�+��{�#���I(@-r��ȒV��M���DǨQ�*��Œ��M��O<&0��w���2�b����y���'�E�;{+������I<��B���O�z��������ej՞&x��@�W��z�ִK��_w�[k�[�C�~��6y|2�2�Db��5G��[���U5��py�dn����Q��٧m�"�4��`�ֆ^+�˙=?��ׇT)���'! ��~ �n�*�uoĕ=�qZ�]�;י��$�\*���>x�D������S^�4����+���{Q�!��?�v�w����r�F:������8*��N�E�­7{�4 ]U�d���h@�&�������_�w�%�mvmX���e��y����l&�x�r��WA��l��ӓ����ZU� ���;�*�FbP�]�{z(O�X�:��4J�z���xa��t��D�Fo�X�a�q~��)�y�ϲ�y�JR�|7`7ã0|֊ex*���v��Bp��,�U�Zm�a�VF�{��&�.NF�������Q���f�>��U��&�Trw�lC�c�Ș��5W�c�]2y\6Uߕ�q�������<�/�U�l�CA��������x%��}���ݵ��s~*�y(��̨il\��������\��p��}��zs$���o��"���������͍ $�J���J��y�E�W=���ǋ��(�5m�y�H�^�	Bt�k���ZK���X(&��M�|�LM���&0��c-uT�j��k[�X�
g��Y�PrW9͌<G�����C�_�f)�ZJ%��ne]�9	9�zO��Ѕ�g��#���� #��UD��Ɓ͐=�@��1���o��f�U�ٜ`/�
�[��nD#����csN5�����(_�~�k7�q���{H)$�s��_3�/��yA�ڹ��s7G�����y��t�`g��Y!�߾���pӝ9G� �d���m����P�X_&��Ok���L�A"�L��2��?q�Cv`0fo`�a羻���iתM0,ia���._�9أ�H�ko3��}���t<�,'��)��mj�>�p>�HC�v�A͉j�τȖ+s;]������*$���[#{e���w整̭��[�[3�G����J��>�Z��E�YӜ}Lp���s�(��RB�� U~���
��&�BZ6s11qh��D���N��\>5k:�Rt�~�Y޵��Zb��rl�ri�<�!���I������
�=���E��*-L����&�����炣���#�|����+�Pk>�b2/���F���`�������]�jt�a��ݎ����g�Y&�So!��1�M������>��3��V��+����d��꿐�����i����
�uN[�g�{*�2Y�^�)L��C�y	����������(��5s�*��)�9&n؈���]�C�QG�A$ЗiK[=-@�8�?q�9�\��a�����Q�(`�����Y���|/�:"˳a�(b���_�����H���I�3�����c*߾IbA�;����l�H���bC�����+�wm%g�wBif�}}� ��5�����Z�G���P "�*�������l!���4 ��qw�|�RGc�O/�ӢwJ��.ŵ9���V���f�H�����?�={��[�9e�q�x��ɯf#B��ẍ�q0�s�^Skr�� �:�t
��ge��`c���55�(��n_�gk��s����v�kf���ǘ�re�}�H`<{1���o
�b2�j;J۲{��J�!Z�o�O�4�j����7z���;[y���L�&U�h�U�����~8����0`����:M[���e0DL���i�.�Wzp!���6|�3�9Dӽ:v��Z�\��˿x+���~(�0~��Ҿ��e�5��K������\��l`cG^cէW��wb�����h��|e�k�k�2�����󘫶�Ă��ZY�[�|��O�*�1�k���7x0���(�4��t-`����'Q�g���+]��%ǌ���� �G��,a�Ɍk?J����y��gis�y��y��d���>��+�ϋ�´��wB���""�r��&ħ�����d��"ᥒ6j��m�[�70�����K�:�UoP����s��X!�)�I��rr|��+J�/�@N��_�2�,���l��)M��f�O��t*�ϭXn>f��|Q����4���J��p�.��w���+>�ϛ>R�`ZW���e�%y79����}R�?��1��ۉ[��WĻ�Q7=��6�rx���ۢ�o-��c�)$��q~��7X"� �VbѫeI�x��J�>�c�;��s|�7eb�5~DR��๴�+5�h��;.�X����(Z�4�2�Yll�3 A�D�q�r��6����G@ 
�,=1&�4h�����~K]��l�٫ւ ��7Xo��uOuZ	�W��n��h��-l�}��i�������^>1���9�%"-~���r�'�"�n7S�ȝ���ٌY�\lF�tq
�U�cӲ�I7�9-�t�~m����\
���f���b�E�����Ɋ���:�^�����(p�J�����}_��fa�>� � ���O���Ŕe��L|����
�2׉���ѠN�\D�~�>Ǆ������f��!:�8���iaķ:�Eϐ2��_3Y�1��s���X�\�~S7#   �����[������-��&涢����{3	�GG-��2i��<A�d�
�������~����ɋ\ ?l@���������X�TV��>s<l��/ڴ񲾣��U�9۶�{n�vE�k^��0�'��[b���T�=�tI_W�'}�X=N���I8m;���m���ڮ���fzTb�'��L8JN�Π_\F��:l�ax�t��5�7�2oݣ[��� d�/*-y�������Z�2���o�:�OA�!�+��f������17e�u_�4(ci��3�'q.*���݊��5"���O�]dt��Eb��Q���D�kQɒg!���FVf��<A������:u��o��u����)��!㮠��IÐ��;��u��զ��ŉ�E2O�H���4G����ˋx�f���{��+G0$�x���L2�`"v�I=�JH���|+~E ��m�.4�ׇy?uП��t���0 ߕ����������-<>G���"�5p���b�h�k���\�_;�_�U���2���7��Os�áD7\�W�]��{�9�R�~{d$�D<��^�ݘ`�p`���a�rP?#���I��E��D�@��ߤ��M{���췡=T��h��'
����P�GeB�؆�Y*=D�gPR}~�8u��A�9V��Qf�����r�j-�=i�5��;~�L��l��LXo��u,j�5;���@�`�YU��#�οr��D��|Y�}_��k&r���������ľ^)Z������~|r�I/gu�����C!�e�ǧ��1A��R�FO�Bu]m�~^	���b�)Ö�ﬔ/�w�X�
�/��o�a�)7��e�)D��O�_���;�:Cw���z�*�>D�m���r8Y�MԺ߬K�1�}W2�`v)Zt���Ȑ���i�s�X!mK���R�r@@�eb�yW�8��h���k��A�ܖ�n��,�I�=J�,����=��O�D?��o��e׊�����9�̗�M�`e��E4�}�Ⱥ�����И]>��aV. ����<���wc����NvXv���>��j��w��W�:O���3���d�u�7S*��h�8�f��ٔ�'�V�fӲ`����aS�e\�W`�&{8�i���ljV^�<x�p��T���EΈ�o���	���X�U]��h\�V�;�0-��'F�����b>�6��KwO���� �d�v� �xC1��Ib������'=��E� �������os���'?p��_|���ejLp#�f|���CE�*.R���S!#�'�$Yy��z�sf�4���ZM��V�u�Bt
D`��0o�g�U�L��vP�-���l��qסh7���إǡ���ŧ�)����s�q s�ϖ���=[^/�\d_���ud�L_a#�jh�/�'m��h��T'guM-��1�v�O��!��캉'�	gz9����lH	����/f4�N� Kۖ��Py�.�u�~���u֡`:�;���ێ�9m����c���[�!K���,(=��,��Hҕ�b�[����D�6�+9\B�8?�]F1��3�d��P��ѐ�r�}A��X����i�-K����Ѱz��x���Q����w�Ϯ8��ܒǩ��۝['Jv�)���pdt�~�ff����6��� x7�鸢d�W��w��!���� Q�"mfwH�B��6j�=�Y+�N�"����٨<��<Ѧ����"��Oq�J�jT�LwD�p�n:��*�����Xt�y�w?C��5!"����� DY4����k�����ʹ����VȔ�iN�Z����������'*����Y����q	��}������j�h�xw�|Y���jb�8R"%l,�S���(/��#O[n|)���ui�����%d�s���et��/88iO�:���X�ۈZ��J��b�
�>�T6ϯd��Z��aB�]��l,q���6�U��5�|����3�:N�W̘�����\��6��O�V�3B_���UA�L��Z��E����ٶR�%��=�mpg�)�)D6&x*�)�T��~ؿ�<���Zl� QI�.��źF��!5����6 �mN�~<��k�Hp�x�f]g.�N{�y��j�>��*���zP������P1��ƝXO�ª���.9���fJ��aK�h�D��6�@��D��q��vS��9�]K>z�3���V�72[��?��:�%���Y�6��DVa*���yP��%��"~/�H����:����33�5�&j^e�bPf4Q���jiX %��Ոz��<�y��P;R�[�x��Z�m��a�Hk�a�"��XO�Q�7���T������O�\�5ฏ$���CS��t�8i"�K�-q#/�.��.�G�+�����iP#�w��.2|Y��=�(_c~4g���T��C�긨���_,VQ��c�Y[�?�h
��z}xC����⃡�*��h�dZJ�\����5�B���vݭ���{�+DD{��9�g��фN��o��!�=#+G#\Ӑ+:��]�x�B�T��vp��)Ӄ��b�z�/����u�[6=B���R���YP�E��=W�yZvd�?2(�賳���p��f]�͔p+Ydj���b�%�^�?F�c��6{�kx�Jڢ*�Vf�k��<b� jG����&�{PUT$�z���-$v|?� �v)�b�oind�~է���/��Gz��Xf�Qe�(Мy�y��_�2�*���	��5t��������^25��T:}�r�ɽx(�2��=y�/{��|��[�j�F����MY� ve�r��LK՝>�m���{Q�_!�)�릱p4h���Yk�O}(�xp}Ļ�p��Vo����c����#\4�����/���>��fnf�c��!q~=gJNp�l�� ��3<_��P�I��rz�[	Id!�n�:n��|����n�%s>;eH������Dn�@7�u/=�;��L��6���j�)� n���Z��|м�Iw�Jղ��b��~a�񳹻Eu��5^jp��,'�%��r��f���z>����g���9�W�n�E#���?I�NXzY����x�x"��.Q^g��u����-�qb�U�>쪤��Ӑ~K{���K�%��}��<^2@I�K��wX��I�3�m�VGa�u �9���e�6V��E,�ġ\D�g���Y�(��ZלI�%�+�-�{Df�*{	�H�W(Naz.P��EyH��GE�"WZ�!�H~C^:��[{���Q����ޜn`zC�B��a����
������6]^U�,?��s��3����hz�}����á�a�ߕmZ'��O؞}�kG�G�G�6`1T������dǓ.�!��~�G�mz�'ӯ�l�bY�<Ў���=�;fݸb�l�º}^[/���4!>�������J�ċ��f�v�ha����0w=������N�~���d���>Rd�*��(�����
��2���wM�7ܓ��ov&Z��m���C���'8�c�c��/��%?�֮���5"����8��'S幦s��T���~�1���/��{>����'�c�^ܮ�����+g�zi���!���jܖg��(���q&4��1������9զRyk�B�d��s�� �yt����g��CTl-'��;>��u!x{P[�?�uq���B��f���1 �ɗ���{��Z�&J�����|�u�D����LI(VOدq�hG�0D�3	��9��C:^Y^)������M�!m�:��$��${a6��AUS� �����Į�|�PE�I�U�b �����M��)N,84�\�����D��7]A����/�8�� ;�.�ϫ#��"ғi�"�>-yr�o�� F����Q�"��G-K_�y�*�)�Q�yΛ��iS0(����T�4�j7�Xih��\�D��jt�ݲ����=l�F�T��)�W��=�ܢd���|�-{1JV�*�yU���ڒ2�Z��������{G���Ϧ�4�А�P�׭���M�Ǚ��ySǙ�T1��_3���Ռ��B!щ�=����ΊQզ��zb*
��k\�h��?d9$*�Va��b���b\�s�J��ً�S��R�L�ZrJ\���s���8�m�@$g����:o�B���4!Ŏ�4�m��`�����4���FL�g���e��Z�\~��l;��sw)����v����3[����L�do�6"�_�3��]�!m&x@�������P�s�b��r�ͮ��C��g�櫎#RÇ.�?��e�{^��ŉW��˥�sz�Ït��;���و
h��p�=�����VH��M�Ϳs��귯���۰VV;��-�3������{�Ő�(��~A~�u��-�:�
��r@E�5�g=+�*{�0��m��r@3��8�d�Ը-��W�4D�rG�[e��uh�����7��F��x
���M��4� ���?�E�L�N�J�Q�6[I�IQ�(X,�kɏw
�>1%������e�'���c�l.pIt���]@�
w�<<(��i����(bI7���SҺ;c��ݺ�]kƇ.&�xE�[�gTK������Ҟs>�d��j� ݮ����Bobb�gg��!W#��a�
��|zc"ѥs�P��طT�̉l���L�8�ʾ��$n�]>2W��'�QBA�(H��ӆ�ͨ��3��;/#��-�bCDؔܟ{�g7��z�U��'�$�c~b��=���<y�F�[~��:_b[�`R-��/����'��=�3(>;�U�A���~��{�o�z��W)+\��n�����Sص��4H�>��R�DR_�]YY4�̀�����tڻ��7��o��P�$�9:F
$�_;i%���E~wR��g5C������Nƹ�/�%�^�L�̳j���^Ň��OΦ��-k�@P*�U�4��l)��ġ�7���Y�Y�����.'n��ո�~O� 9 C8v���fvoW6ŧ�����<���n�!�$��sr�l���5�t����h�bG��4��\�^����輌*���e���q�
#��8�)�����lQqS �r�Lv3��D�Y*>�v��e\̤�\��{�6�|��P����|��NI�XTS`���5�|̡Ll��4��e�CX��c~%�_�e�r"Vi$/4�k�l��s}����qH�jQX�D�0��>�F�Ƿ�F30^����H�r�m�ҏ�������e�mSX[���#��h�Z6g�VĽi��B����z-kt��&��e9F����LVno�l��yB�����W��^/X�>[1��O;DI�&��n��D��@5o�W��룺z}�8t�<���g��w��������u�>��tx�OH�ZD����}�gyy��Q:S�b`Sn�3�3�(ާ��=���/�v+�;�9
��AI׈_���V��c��QZs�Ӗ`,��
~7��0�����sV0;��L2�n���pː@�5;wBKK}�@�����P+9�6���ә>��6O�{�U��BH:ժW��$�ڠi�"�@]�lx~������'�;�e�~�*�4�<d�}�R3��R�qD�E$��K�Ad��,�^)E�a���jo�q�3�E�XW޸uP�.�@�k�a��0r��|�����.�=�ZD��=!}�T�M�F1]D���Z��w_�}����^����4m&��̂�0�g�oF���y%h}��@�.v!P3��/f��yg;��$J�6�6pQ�9״�����koi����B����5�>�u'�V�K=?=��~0Xf�+��uG���:c�'��D�[��7�_�/�+nqn�	n
��:+��"/-� �{ǽ8�?��=�ɭD�Ƅ P�x��aG�Im��u��~}vq�2�7��]����$�����N�����#_�a
/H�j����y7�/�En;kOD-Q�<L.����^���NV��Ë���E([�Ύz�Yؗ\A�H���cґ>��Y��M��Ob��V��Y�'''Y��y�%�ư0��JIQmq+F�� #�O���Q��r�@~�H(�H7�v�"�IՏttXc8H	8�6�gb#s1�b{��^��Yj���2�=�+���̸
�Bj��e<YQ�sWeh7�(1������Q��j�sUԠ5�
��2躇CD��wL2�!�L�k��)�j�5��POȳF�Z<_xA7t�=X�;�궍��`��Օ)꽦�׹�ϛ ����ԫ��ɌY��gm��\Ջ���Z�p]xE\���ް�Z3@�ݳ�Ã1��%�	7V�4�%�+�(���6z���&�N!��9��ܑj�;�e�tG���1���?�L�mBRx��?˅��'ze��%D"�bY�.Pͳ�s��y���7���j�y4�u��1Ր��VU��>��!�7��\���C#�S ,ַd���
��M�l������U�"(�t��|���˵�B\z��Gt�������d'+�y����~u͞ �������}�C��އ{ҕ���K3�"��&6�>�]/�"� �^����#H����v⤘�h4v��F��S�� ��ONXN�tx�~������d!X���o.�ʰ߁�r����v�n*h���=��u�aT��6�Pk�FKK[e:�u1|���h�ݷF.SLu�Y8��M�njJ�9�W.��"O�P�ɚ�k���z�Y%�B��1=�Ma]Lۊ(A�QwJ�&��Y[I-2" �ޟ�I�^�~2χ��Co����+W��[x'^�J~I�R���>���u}�u�C]$ȹ�H9��]�䂟TC4� _�1f�%*�}��<k\�3$�����
_s&�B�r(1V�C���5�:@�?��V|D�۰�e��3Cč���L #+Y9��g�F���1ǥ8ǣ��}Z.�X�oL;��ᎎ=F �Oϵ|����MǙG~ϑ��J�e�M���Ñ��eۘ0\���
��^��˷�X���QM���d�����nvw���/�7ރ쁖�����Gy2h���K�1 w��t�耸d%f£��ׁ����j7^.2�̈́��\���_�d����9l}�?�2�#|)�|��������B���,I�� �s���ՀX�Q��*����}�~n\<�F�0���x��3��y�ke�=g/{\	*w�+���k��ѫ�u[�fOV.�ө}x�?prf���Yt���p���!�[��Vq�3,�' @�쇉�e��ٵ�#��mO#dgJ4�Z�)[����-�C�Vr��rF�N9js]5ng)�R#�>��1����zU?Tޜu�{w2p2.�k����v�lקR�U�- 5Β@�����իs��ҁ�*�I��"�a��p�@���`PC2i|@����<7R�j���k�ᘱ.]����Wȅ[ (�\}��z�����X�I���0�*:5	�cy��9�
���2h����oS�`T�	�+>�ڈ:�Y�?<|�ŉ��R�g�.���g�$$���e�ޡ�egli��n*{[W>��C�;=.nf�����������6��~��.��(�OQL��]dU�>7�H�
�dE(�r 1o6>��Q�ё;!A���~���k\�s���̊���Z�������p���~�Cuy9R��D>2�<�ejf����:zg遃fS���pAr���Ez��9�ް�&Њ��T9c"�A:ǒ�|�܃�!�"�mW$U��.s��a�XR�?�Y��Qn�����V�0N����?��p�a{�h]��'@��ODH���T�3��x�:F�66��r���\m�w�[,�aC�o���(v(=� � 8����V����x�BY��OF�4��~�V��� ۓ����y��QO��[�+;UWo3n>��@:�kJ��3���!��!ϸ���z�>�{�(�����< y+i�F�*<"�]T�0b�#��9tN��X�òN��E���.��d����~�0���V�t(����(L_�y)#��]��� ��䯃�ӡ.$�q4&G]�'�"����x��@�M��}$�t��hy+���O���(J:dR~[�T�ԋ��~Vs�Z�~`b���^t6��̽�L��mƇL2�O���V/���^]w��C&�	�}�YP�kc��Z��`w��5�Ӎ�¨�sBF͊ޱL�[�\K�����@D�J-���x�zˌ��d���y�i'����ղ#h!���N�<���a���ȿ���3�,|c/5��[�k��&݉)����}����!��Aĸ����=x����R̹ɻ�?�~N�B�U�eB~e�������;:z�U�O��_��(�JB���%!e��v����5*�̤�W�W�y�d]�Y׺6׺�v�������~��z��|>�9�׫��=�Nj ���:����E[�33w�m-��?��㉼�肬-]"Hg��(��M�o}��.��Ǒ��VZ�Dg�JZ��~)U��Q���Xh���Ƈ���65	x��1ۮ6F��)	#�K�?{�����ZI�bR`�ˠ烼�0V<�����j�$��r�eV���ӣ^�ߤK�z{ϲ�n��R女8z^nZ��$.ö`T����i	�[�����>�5B3��+�{�:�֔�q�;��,�J�=��W���Pw7ָ%�_ �xe�9�:�8��V1S;�����aW(+bX ]�&e�EsU���㶩.����4�V��h3g�0�=+r]�&�����j#����D�=]}	�mFȁ�z#��ف*��f)�R8Q=�V�=Y©:*]y˓�/ls?,X�r�$JZv�U/�;��t���i��A�����aW�����I� o�q��(��`Yd@_$�%jvzW��HP<2�LY�c+kWX�f���`s>�Cl?\l>��:)`�._U���x�2z�G��)�1>��(�vwT����˅�45~���͜e�a��~!�37ނ~��p�/o��R��j[�8�)�.��18����0#��̩h��ɵ^�J{5C�mώ�"猃y��	+H��jp�Eǜ'n�b �E�4? �=suRt�5
�D�ѝ����9�g~7:j�4��������W���l傭P��Cң#�*n�`�4�ŕZ��C Pa1��
���k&�r�f�d��a�W�芃�^�O��V�pڼ²���HƳ�hL=�0~o���4��Ꙣ�̎���s7i�!O�?�P�qp3��-�.j�jH������._���n��¤�_�~~`�17a<��[�A>l\�؜���ޏ�r�����uP+u�|̏1^_���weQZ����Y�݈%p����j�p >9�`9��� H5���6e�G���R^�7qWn��1�����mf�2}�Fmߑ��{C	h�L鎯��&9����H��t"�D����ƃ���X[���]Sz�!1ǐ��AJ9%s�ѸzjA/E"jܣsw�&��%�g����Wn����S �D��J����4����j�:�Z��w�z�.�\tUM��y��#��4��*�uX^lY�Î���r�7�����l}UK�����w:�˻�����O�,t>���K�����/l�]�6�Z���>P_3~H��gO�;���A	8;1)^�J���؄#0��ߜD���
o��Z�#�g�r�Ȃ�+,7��2�K堕���Å/]�����h^f���}�w�t�\���r����!v�.h_�]>������	=����e����OO�Y��Őݮ�����ݗŉ���Y7G��oG�&=�먒=3vN�l����f�W�KߏէA�P�i�f���	?�M�?��:X��
��JZz�eJ-�Ek��:��3t�,!
�]s��{��w��YlL� ����.k�L���1�w��vGz�$x�R�kt5�{�"��D�4�l���_�ߗ�,����xR/�8���֌��	�وˍ����x�>����[P�5���gU޵����uT&�T7�M������ț���@�eiϰCso�A7��, p&��i�9$� �d-V�A��xTV��G2�+rZ�
��g	ڷz��4��1ݺ�$U�})E�"��J�ġ(s`�����(?\m��˰DJ�}�/�}��'3rh9���������Sm[�R=�Ԧ#����j�v(yw�4�� O�lԠ�h��1�b>��>LSՃE��I��r���5��l?�F���P����W[��i
_��P�i�e�����sG
hF2���,n͞�~P���E�>�qe1#q&�z�;}��_��� &�8�,ܘ��:.��eQ��.O�������u5������6V:�g�4�8�L�SE���s|]�b���3�/h���6�s$�kd�R�����!�h�s�1<��ay�#�B5�i��A���} YE�dhfnO��$��^o��*+�Kv+f���h�K�&;v7	�r�ý�#$�� ݷƯY���ߊH��lb�bՆ�=ia��1Rf��T�!���Uo}��T�-sv�N?�b�Yn�d��T}���K�c�ч�v^�2�KՔ��O���V��-x�#�U���W@B�5��g����=R���o��w�N�I������q�z�c2���}&c݁�5M���]���ćR����5�s}T}��Fit:�^ U��Q�#�T���r�w�;�|���]��ت�4�R���Suz�5t�8�)�{����1{&�e�m���ҡZ�̳��QX?Z��:�<d��~gj#����5���tۋ��X�ޯ�
Q0�kS�m;�nۥ�^4��}��G�}$w����f��t��w�x���mB��viF��vGщZ���.Db�H��Oh8�ܾX'���3�1Ӝ���\���B��	nn���	���Awën���)�A�b.�=xi���Umm!��k��¸�[s������E�3����7$N-!��Z"i�Ux�B�-���������ǀOh���G�.�J@f��N�K����j�c������w�C	s����c����3�3GK�X�*���m�^���e�>�� ]p�zA~��mO4V���2+�zŰ[׼_���tܦ��O�㾥��)�<�PM�yV9�!'~)�{������_��%ݩ��wo���s�42`	$��?�9���0Fx��𭌳c8b��З�6ɠO��y��h�ϽfҰ �'1GfKݺ� ���az��\�WM*Po��)/x��fP׽ ��Ѫ�w��;��Ƽ�W%��Cz��%O2Ϭ���{I���s��T��#��e�NB>M����ȯ����I��R���׋��i
xF;$`�~|ے�T�L/�Y]��C{AQ�e�Ü��7jN�uW3-Z�2�-�;�"����s)dyP�=�2÷�������Q������)G`*�X�T-o����՝Պ��NS���b�q��x���Y�ц��/�7oh�Aτ+�@z�A=/{�y@H���g(
����`�o9���hw�l�Gҋ/H/�������.h�]j�='�>O��g�j�%a�̺�����~8�q��WK��Ю���`]ܤ��ccΩMG��[T1s�LZ\�5�����#�1���.'����g��&�9���A�Z���'�a�f�q��F[�A7�j�ͣ�5HD�뾄�'D� 94������Y��;XI�&��Od.8ʄJ�ӛ[�-�3�\���}2�-Tc�Y~K����32�1B%q�O��I��u��yƹ.�Ǿ<r�����-�8L�����3�f��o~,O�i_�]���Ҕ�4�d� E�����^��m����HB������^��%�.�F����%�B}{
s���VD����[�V�!N�6ƫ\�8���#OG�޷�
Ӳ=L���jo� ��z=
��9�������]�_����^��������kƺ���y�o����I $O�OE]��{L�<|��|�w�����QH@~Q��X�a�͈��?���6�_�����"��l�2^�?�Kc�XK���n.nZ>���:���E�p�1f�3�o9� ��3ur6}8)�&k�\#�m�����&-�kv�a�X�uL���1IaC�����gR7�4�+:9������m����ZF�������Ξ��W�腭�,ӲP�1<�#��U>�q��5�BL�kʲ���ݫ����cd�B{�r�tm���\���)?��bY$��a�_"��hG�	��v`�&����Ok�;���{�B/�����6��f�\�l��E�wl�cF���-������QI�iu�%���U��ٞg���ә���*�UD(L3��C!X6`�]�A�y7_ߏN�Y�Ќh��f]w	B���nC�n�}�;�C�HAD��a�K~�Q,%�9�Mꚿ���70h&m��\H]����/���	K�13MX�n|@lL(N��^e U�R9�����^>�b.�&��S�y�~�Ru�:�
��6�R�
���(���-�^�ρ�m ��G�:Ps��7;���w`� ��qs��Mg��/���56&OF�:�V��C�i�W�%��i�O�����OjM�#ge��i�����f��Vy�Eh�K�i�
�ae搤�V_<���&��.���F�m3� �3�M�I}���� ��":U�g�eR�_kc>Nk���9��6��S�n��D܍\��o�?����"��?R\+�2߬ۓXKnnq���v��N��oL\h��b���KX�L�-�V��,M��x��/V�.�=�~�Igݰ�c�����CH����1�ͼ���L��������7�����Z8`R>�:aG�h�8R��&�Y�[V���XoP�3Ѧ���rn4@���C-j��`���j�z	rDO�0�d+�Gs���\���D�Xos�k�n�5(� 05�j�+n�~���V1�=:�۫w�X!2|OX�U�҃k�z�b#į�mTJ��|7��U���j?���^����m�a,=�Q����o����6xπ��y�d��n����U�Qh�庚c�r�z�.9UH����ڢ�|)��m�B�4=�^��m�&\a᛬�b4%��'2��� ����t�v_笻�Jg����B��<d�]�c�K�Y<Ig��e��rp�'��h� FH�tC�{S,n��LqPfRƂ�-��ww:��,��:��,�sg<_W����4H#���t‶i�� �p�e��P
Ou���s�O�RFY��M����t:��,�V�5alޅp�j530��U�cRi�\���>��5�>���;�U`����x�ܨ�~x�>����	�m��&�O�y,t�FIX� ��%z���Ү�|���2~�tا�ȷ>y����~o�4��u?|��Uj�#^4.�R�w�X�]a'8�sA�����7��#�����g�ո��:>
�"ptY͞���ya���!K��$���W��)I�ݼ���>�B�PDɦ�� ��FSMM�"X`$7fey��p�m(�ѧ�Paپ��|�^�p���9qo���oa4���J�r��Y�V�-�M9Qǜp&�t��|�\g<G�ā
�.1�RP����b�TS]N���=N�d1C����>v+�z&2�q�i¡��=FL&T�t|8N�S^�:K���A����e+�W���@�3V�>�ʹ���S1��V^�&�fu�ݤ��SJRD��N���`�@���-"�o�M��g�=��d�<l�	R��Zc�u{����En3��պP�@����~`L�M�U�S�p���n�=�ǤD"�U� �@�O�X_��Ń�KoG'�GO�����6�ˇ#g�\0���h�[���ҋI�]�p>~wZ �����4x�v�5���ZD�a��UC�{�E*��K�<�z��8�4��x�p�E5��֒��S�k�������	N�;����kKq3��I��W�c��D��π,=:���3�J0N�Q�GV�R�)h0O�G�R�����f��ޅ�6�@��mO���u��Ɓ}J��N6����Ό�_�7�u�k���?>��ho��L����nvL�[n�Z9\�S�����<�@n���f�)�N���	W�gقR��������?��=ȓ�P�.u�SŒ �+=@c���@��2�q1��82�~��>�l�b2����{��<�kY��e�tܫ�n�#_�P,t�m����ba<���Ą��	�|�Qtu���-t�W���*�O���h�LB���~J2!w��35��ձ���hm6�f
�`����伺�mQk�{t�y����Rяh�.����!����M�D��(��E�|�/#2�|�>
KG�{��N�5\�ݾ�T��QR[�I���=R��^#t!R�,;K����9�֣z�. Hm�
�͸�b1��(L�Pe�t���*{O$�rXۙqT[���2g���vCy%g1Ә�6���p��#?������o�>��L���oi(�R���):�J}Xbk�o�A�+A��P��#��������oV���"ĵ�2�*��e�l��6���v�ؙ�B.��x;^OH� �{OG+��i�FO��@}��ow����j�x��y9^�I��le������I���E�D'�S`[��<�D:���H1Ы��	-���e������J�j���wp����okFM�A��D_�[����9R<� ��"Cu{�
��D�	��S"4�+Dqp�6|��Y2Eep�/9�M�"��+��ky�+I�?��%r�B7�ȶG~�)��\v��l��pn���m�Z3��xi0 ���x���\���DJJ.s���~;�w��I'~���]��j���>���5z�A��$����0�_I�����ʫ��1q�w�����\"_���̫F[-K/n������\z��P����ܶ�_ϗ������at3��AR�Ej>+��DA��G�n�������]�ð 9t�A��z7f%�|�<���Eq�e��i���D���Z��E�J����lm��脸0���孆�\��^G��
"b�i���'�E��%Ao��&�o_��x����}��$ak�\r��h��K��+�q��¨C�?�ʯi&�bV�Qm�0���9 ���K��0`?��.9��>��o�C?��b�~X�h�{gt�JD��%踯m��)�]��
�˖\�D)u݅"�\��I�G]�8����ǂ{w��ya�ih�d�#�5�j_��=SkUԭ,�#$�[�(x��Cq|��*uqBF�s���w�t�od�c&$2͇M�`q�oE��pʕ��G嬍�ߍ��G����Oԣhx��+^Y��\L'|�Q�P^8+�U������P���)۸'2��p=^��^I)�7��Ђ��Bi{��J.9�Ű�
-�aqS9[�� 0{��ש6| �s|�tl����*�J7��@4/{���I[u��6��Z���ʎ�|Q0&��Gx_�c�7q��SG�R�s#�ɢ��(H�o	CK3o�U/է7��Dm��if�A`y�@��(~�q&��DL�Ejg7��vz�q5��� 6g�X6yp��4�\^��u�NW�Vd�kd��$�|E�+�L�AL��˃01�aд�Ҳ1�dsq
o�]��?'._5��pgqa��:h  �����%�aɱ.G��6�v��VVp^l�g]Y�O9f�vno��C����L������%��$�]�l�ܨ���a��-��kK�i�c_@��B�u_�����/u���]��<�XE�1������:�oָ��Su	������܇��D����+�/���y���\w<޸��KPyX撼��̩2�C��8�<���O��l��R���K�,���"��B����{�����R�V.-5K��h�����
~��椩�����08�x��~����у�sCȟIym0��tQ��$�*�y��Λ��)��E�N��B���)����ɺ��[3��N�� ���lQO�:I��q\�io/u5����P���t�'Yq�adw�Nx���:8`O��#mA����=������e'5e�x��
`��@rH>��	��d�4>�ƝN������_�&�٭+K�����W�hvy�<ǝ��c�gvY�;prr4��vYt��;�J��6H
�.�Խ��l	#�v`X��?�R�6�[�)5��MUps�.G��"�\��9L�R������-W�~ܒw�C�I�`s`�����%�ؙ�&R��#;���'�sj�g@C�_ ���s��C�4cs�$�F��z#g�N7��dyOk���n6�Z�]Ϥ$|���>�k�2�z���
��m���5����#^4� IR
�iX�k���W����R2���J9Fo�RCc�G�u���lH��[t�#�D������}����4�X�)���n!@Wv�I�	F���ރ���9�5���S^R��֧|4��'?"RA?��.x�1��Avu��������+.S���;K�_*�j�[�@�c<��}Ͻ%G*���R�J���jĢ�i��Ko��6��OcΫ/�%�*�9��|�.t��N����,�8�~[��\�r��ů��	�O@��b��u��J��4o{�!�1��c�1�����\������۫�n��\r�R�#�π�
S�����s+��͟��1�/�vg��iFeB9����!���_���oI�����>�R��{&��Un��� {V]qYW��0��2aj���<�{�H���a�|�ӱ���JN
��d��bi�B�oËx׽��2����Pٷm��b���s�ue$Dç�`�瀭�E���fT���0�SHJ뚢��*��<��-����*�p���|��ፂ�x\$�u!�X���z��>�a�!ƥ��#5�7J��i���jur�(��Ҡ�����(���lg�W�c��W�Dݾ5�F������,ԊP~!���(�����d�s"����[z��_��_���Di�m]^ֶ�l���~��~�}'`���|�2ڧJ�@�������4�Nݮ�O��`V:{H��n&X¹1��:��0%s4
��?�'u@Q�A�� G))y�enԸB�L��fl��J\�e׃��<*+y1��Os�Q��<��\��{l�/s��sO��JP�կ|AK��x�
���Pn�=���d�J����ݖ�x�a�x��.� ���%��y�d�)�Z�ָa1���,�]�L��1�K�O�o��Oc������8OYjY�GЬ�,E����Cڄ+,�����Р�MQ�f���Zߣ��~]>�9o9���>pջ�p��r�ڿ�v�' j�cF���H���~��n���9A޸�j����_3����l�C�!<'	G�ӗh������P�P4NS`�mו����w����Qp��xMJY�	�������ێ6ho�ֶ���,%n��v�nk>��?�$��h���x^ �AD��7/K���<��m�^�J�������[B��K���,�t��}��^�I8�H_��k%�����u+����|�����#�m�DF[�'��܏[�c��OӇ>^������u�$�X(�m%�أ1Tu����˅o�ly�߫ȯ��IB3dH쬯O[�H�a�n���>������;�!~O��m�_�Z�\����Mö%�x8����/��DV`�w��1��1j����5_~�|����t��R���"vn�p?���Jbr_���=���r	�_�{*�A��,	HO��|Z��=���B�[|�d۠��5"Ӥ�X�Z��	�zu���W�W��ð�斿B�;�R�>BLW5	�����{<K0��H+O��<���,c�m��u������kE�U�)/��N�D	��Ox^ã`����TS�~ɍ��#5��2�~����k=�&gB3X�i�:�Ҽ0\m�3C�r�4`���Eһ��R6g��	�	�t�]���Q�A��吿���vvM>��cd(���ˤ\KM�ٟ	��?�O�Դ_�t��i��V�9��e����õ����9?,���w�/}� O�8��*��[�&;;�9A&���t��!��|N΅�3^r*c =�}<�ջ�'����e�^uG�V�Տ�.�C���l���ov��z���Ѝ�B���^�W�Dl��CL�ky���19_���t�Ȃ55����y��CHC#Ȋ���s�\��Z�y �����i��|���������K!0A�_���B_������#Y���%'@?�J��hu|R\zl��J���?�Ɉ�2p�~��#��dop_�)J�ܾ�V>��iA
he���_�����R~~2��	.��K~#_b���=:��/��Z�݇A��@�/&#	ǥ�<�Q �O^U1��O����w+OZn,Q��xLà�C�}Ӗm�}��Pb�3�4�K6�Wf9L��	o>��D8�CC}�F��eO��"�������R&�e7l��=��QU��u�R�@۾O�L� d8�l�պ}!K�.ǂ`7�s	��1X��ORZo��ղ�ba�عn�Z��P;<P#5�$Q���u���d�Dx1P2K� �]"�}�V'�W�l9�n�+�|<Eߺ�|�D�13rp|��$�Ts�2Z�ܔU����i�g�Х�x�;٪�}7v-@?�ڌ�wm��a�$�ٜ��e��SL�s��ⴋ�u�����ӺOѼ�s��?iL��8�?�h5o<�B��[}��d�z���ܹk�M��J�[fj�!�U���d2����IY?e�hZ���|�� ����gxUh!��g
zq�C3�c,ѽ�Aɳ�R �j{��r�ߐ]����КHs.R�۟���-VZdN��,'���O]���Z��<�����_V^]�����\����M����x��5o��@�1.��ʥX`[��x� w��x�CiRǉ{xn�)��s��w��"�R$x4�¦T���=���j����5.�"L\4�L��ugo�c^S�r;W���&���`�{���=���=�<jQ��JI�ΚJK��1��^���B�&]�O!��3(�Bb�0�k�ؠ��Z���wK_U��G���Fk@��C���u"s(�v�|��js��{�W��'	�XG;Q��*�T����<ƶ+j�>���2���WTV1�[ʕ��U8��Y�.�9 c(����i�uh��������e!�M�Z�G)�����.OE��Hu��N*MEe�`H&��?L6��@x�<��A
i�PA���0��t�/7�J7�_�������hd��4r�1뾅rhF�&�h/�(j��F�S]%4���"���W$�\�_z���)�OCcEHz}��HaF��e�y���ظ��W��4��R&@����iņ@�5�}�_�(�,�j}�Z.g�BżaR�^Gp�x�n|�I"���:�Hj��lU�?D���� �c{gp���]��-�_���Q7����U��ho/.��񬩫�C��<�z�o���ub�y�����>r�t	�no�(�
ϔ�uvv$c1��u'?A�߼�߹�\��}@�l�iy��/xt��[��]J;��>`�:Oy6<�9e��G����N����Hӡ�/�e*�WV�'��e����|Y����+W)L�gXM���+��=�"@m	  �lM!�c�4�`�������)�(�)���&��-��A�F��Ǫ�:Ьw�&��k�?.Qu+6-,�?kɏ���x/��`\��\���vc@�I�>��dp��u}]�H��3:D[L�#ɠA�uLN)��X����B�X%vrs}��%�����ab���0���t�NX�zs���f�f�,O}P��k�T��;d��c����"u+�*��:=��Z��PD�G��w܄�0g�QIH����5�#�s���hl��z�3;x��_���Ѡ"�L����-zc�ʐ���s�cX��q!�H�U(f�xǒ��}�Ou���֮Z�m6H��.8��C��-J�CY�ʟ�������8���߯��lsR�<*;3ٖ���Ϳ��c�~���P�;5����jj��]�k��g��C>R��y3?~v�ǩ�����(&���9S��N��j�BM a!��U'w�h;�cl%�h�"���XVVg֓G�M��4q2��g@����?MAm�4�Fl�j�u�ퟏ��[���JچX��W�z>		�Tx����y���8���w^�m�'nOX�|('%8���&u ��o�&%?\��KRHl�U;3zW/I����K�{��HYd����K�l��:Y�К�_���B}<Ź�A�~�e�1lB�$��nV�"KK&l�3�2���\�L��O�3Z묣��>�}�F��u���l��?NUʬf�K��KBQJ�&��A�1;�M<�����۾�2p�}>��Z$����F&oKo������:o������i�ѿ�8�j`8��{J���o$ҿ���[�抾e��V��$n�6���dM�a��7��σ�9�28/-Z/��d�����T\�&�7���H	)�h��.��U��ǌ�,�x�n����sa���_��ւk~���4�Vzz;�U�۷���+�VVVv���-#b����r}Sdr|��V��4��.��ea��)����vll,M�u�ܕEX�w�*�]rƩ�3���8�X���+�E�| ��ru}+�ˣ*��&W2<1�W�BEnb�9�m�T�B�a	���٘5�Z���R�{�.O��R�FKYE=��}�"s6ZNU�>Ef��7A_!�lִZ�]<*�wi�n�p)���Ci���́ �ֻ{u�,��p�h	�A�}v�4s//�|!6�6���\�K����5�W�e��D
J��_�yU���K}��V���tŵށl��H����(��RȪ_%�<�wN�ڂ��F���Hu�U'0�Ey�S��J�h�ۑͺ]�f���Z�"g�n��M�RT` �x�ܟ^$4��X��4�!��b���`��1��S�/E�h6p�惑.�~�9"�[쾚���P�V�U'<�ŏ���i�>洣���G�(�|�Q�z�3HYX�˕�u���p� �MZ�t5L�Q�=dy��5ߣ5�vjJJ�i�����T���'g#�̡�������Ã�~����yG�����c�o�X�n����.�4�,m���2������;��.�o��(� Z�yin)�l�?����O=I���r�� ��
c �{\���M��%$./�4���y� �0|熕�UsX�����p���%{�e0	H���,���.�pчS��a�ۙ�ء�-�Vm?�N��Z������T#��qЉ/�yUy�gw�ћ*�
����!n�v�gc����x>��"��w$�ߔf_H�o���	7�r\����/.��ow��9<TL�����nE��.|syUMnQ����aw{�q�3�2:��nB.�hz���6�2����fO\�(�#`V�7kd�y��[�D� �B���m����t|y�����>�Pey�W�����.���K����	���;:c��81��7��J��vgC�h��6�w5&���P�|�<��(%�#��G>f5���	4AzV!:����>��{�'ˬ�û׭�k{qu�E�uڐP�%�Z��֦�<�n~����=��9��Ȑ)'�8nh�t�y�&g�,<pvr��Q�)��k7��c���143_n��(n� 	L� ��e�.ˡ��x����q[F=��S�6�i��������~�蒛�h���I�\��h�|���F�@Cf��u������\{�͸SZ��'0|��*bA��.���<��v�D���w- ~��5�,�/F�~e��*�U��2�'ung����@��	�����\������S�.�yH�i���f��M���c�]��0NM��r�fˀ����x����O��3�.F1���)@�����M��u] ƸY��a�
F	��s�_��m�D��V���C���PȥWV�gb7�X>]H�9��`,�A��f�p��'jn/����{'�X9P��~̻h╞/4:�G�K�~u�����_�r����3�3�@��z.�m�+����}U��wǣ���k�Z�Z�cZqZ$�C��+;�I[����7&0k��|��M�.1`���K�?s���Ix3#:�Wlh8�q==r��#����gdE�<�I��H]�ޮ��{.2��̿��ܔQ������D//Q��r��h���U٭5�K9l���(��ʀ�oC�,�e�t��C^�� ;}ğ�GP1���s��ҙ���o�j[�vY�[� �w�䐒�&i|�B�%f��"���B$�K����evҬ)#�1�l�'[C~D
,#�SGK����L=�Ǫ4	o�]�7I���	T���Jc1J0/�J_�k�/�[j"��KEH<`;VH��\�x�Z�3���k�o�݃²���q]8����.���*>x�c�W�J���\K�U���>>�"I�k�5��8�x3q�S��<�w�yG�U���<��;�h�΀f���b�R5n'5���vU�j_CǴ&��G* k1�USA� ��<tdRCnU�s�Ə��L7~O=��Jd���3>#�DU�e��C�O�	4w����̓����c-mu�vF�O������[w:}�#�'� C{�w��	{��RE������ɧ��|0P����8�H�+
J�w���++�s�3��?�矜%i�d<�s�(/:S#�ϟ�
��#�FSty`�"ˎI�s� �R�L��-R� 1 ���,���>
��il���&v?�$E�A���3"��6T�+%V�Ny$�vY�VڷL��`����J4u������eA&�UK�p����h���_�1Z�U�U�����Ǹn�x����c�#t��%��핺&��$[>�o�؉�9�Ы��	k72\�G*���>�1i�ҩQ���Y�S���>�T9U!�� �O�
�����o��H���v�(���"��w{'��}�"�*�^N����$Z�.��#��M����p,�\��X$�Z*�)	�����b�<؂U[R[f���e+&Ak�=e��KL��̉�1Q3��!����]�4��"����A�螢bt�,��Na-Rt<����%ߛ�O��d&?|�U���2�����A3,�"�=�Lt��c�ɐߓ�i0JC2���x/o�q�n↗���0i����R�KE�oߩ67�	!u+�O�t8�Rkq:hޤU�fߪBMR�����!�(�%�id�!&*��>Dqun�	�g�e=�<�{�#t��d�1b�KW�?r?��y���loo��0�+�;��x�NU+3B��많�b�VВ<�/V��ǥv��br��z[���j��;r�L��o�&���Ľ1V��`U�ת��N���{K���3L)>��hsl�4s�/�yȈF���Du+��p�wݸz��3mh����jca�n�3�}���F�֮p�J
?�J�;h���6>Yx--ڬ�6��R�i��*��v��}}2�~O�՗�՗�!��_6��dC�����<?+//�j��IШ���V� 築0�D��K���E���B&�}}���n߅$pq\TF�t�_`rM���$���(#�&���kf�����leB�O�B�P�叭GE�Q�x;�8qΨ�{�q�s�&�W����0�&�&�B�;1{q����T*�@���(��b��]�%��_(�;e��\���&	8Bzem!����_K� ����$5͏m7�:w4枕�C��)B[�:��5�
�9�W�<�J��Rw�.���ʳA؟
J�(|S����>8q��"�xJ��)(�c'�yqxK>W��U�%�H �iܔ^o�.$��`RW'\���R����u���t~D�q5#Ku����Ț�[��j���"�j��)Otrj��h���tf�P�4@�j�����$�1˻Q��p[��e���_��2����OUh�T�����쐐Z�>�8����+�2��R�=x.�,�+��MB��'�������`�Cv{AL&�g��^��3��P�cUP��Q�xI���YP�En<��1�M��Fu� _�%K�w����1��#w�_��C)y�s�ӓuM�ɿ��C�`���H��3�0�l�����Ԋ�����f���uS� ��~ؖ��ؽ�h�'�_��$��?l�A�(lg$�5�j�ݳ��#g6[�'$z�ϯSed�Ӧ�HA���j����S�J�;tK����u�JHe ��zR�I��<���8RfND������De�2̡�S�խ���Z,-�G����
�ؐ���NF�L1|���BT�I�������4�fx>ۙгX�E7��H�p�4;3Q���(^K��pL=qv�g!m���O �������ַ�S��.m�y�����aI��o;.��fGG�d*�N������z�������K��{M��>Ҋa�PF�w�u�xR�ԻEY��s|]��9㭦�h����U�g`I�xnv����C�\�}�.a���4��%�w;�ZW���:Ղm�dؕ�c��'��bg_�	f�I���:�bw)��S��D1��8��M�GapF�ۖi�� :0�仄��ܓL��W��(��]�T���"q�pK�I���gR�tپ\�����g-.����z�xx��4A,LHL|v[�^?��e+��w	�t��yY�W#����q\����\w\	�9��j��fJ�[kߛw[�䐢Т�U��I��j8��,�p<�o�W�?��d��)�J�@�p�����§�mtB��ں�w}���`\�1�|S��}�$�ÁF1J�PQ���	le�7TvY��7L��x-���������A��79���v�A��/��ίS�|��yʢ��69[��xs��0����� � j�E���ѶprY��8\���-�ޖ����P�lyc��ܐ��XRɍ0�}Kqo��SmX0y���M��%����ި���k�cQ��^�ݏQ��Ǻ�-�炲I�t�3�8��U%0������3,->�]0�7>��x������(��--�m���[��6r�ݻ}��6{�(�{ȃ���f}ɯ���<��^.�Wl��?"�=�����;�I*��{I��aT�ʭr�r����F%$���r�Mb��$�un�0��ƌ����7�������<��8��|��K��׻u��_���XO�Y�[zw$�y���+���gևQ=i��{'��y;Y)�ц�������-�����{���I��d����,]2�j��+Y���_��v����W����Y�K�����=��q��?ߞX�F3Y#��wմ&��v�Є�z��4sz��;��<��yLrF�k��M:��`z(Z�����6S��2L�تoϡ���cʟ�������I��1񈎠"��V�T�N]�G���3;�ny>j\�.:����a Y1d<1��#�;:V��u5 ����I��O��"�Gh}J�oo���9�������1<���Ξ�9�c<�*��*Z^�;Y/9�V����,a܍FĆ�Cp��[�X�ʭ����Q�1���<�q�!>�5�$垥�ƨ�-?	�>LQ̓s�b����f�n�﷾�y>�Ǘ��{v���ul��N�V�o�i��q-Fl%Y�~+&7SV/+�B\�[E����^���q|��=q�dݳ���SK�L�������γ}R���tI6��f��b�c0`�I6oH)޷X�1����Ѥ3h\h��B~�POY Y1�o�5�	k��3n7��1`2�lC�f^.i��|�����B�Δ����y��C0��ȓY\���Q�����YK�;��A)���>P܃�y��à���5�z�㼷��_�_����@?q�g��(R�%�5D�)���XA�&]��Y9
 �xe�/?N57^7�j|�qn�n �퉬��7by�兞!�Ϻy�J�[��V�|�N���	B6��+�O���>����.ua�*����I������>VU3ȑ8�����:K�c8}W�ydE�f�n�:�v癤��v�x���}�;6�&(��\�Yޫ�Ϭ���{��y6*� �܉7gyK�[S�k*�!���kg�e�>�<�����k��m�F}�v�I�0�U��&��1Z���;T�R��y�(y7-r�}�&/� ��WS�8���C40�Mv���,zв1�}����M$����VfI�ɽ�Ϭ�LѸO�-]}�X��v�}�dt;��o�**Fqr�W>g�׀�q?e�����ϣ9��|Q��x�ۺZ�}��0��|�:H�X�!����.��De�߄�g����nR��&�ZYD=�c���2yw�cJbgU+����K�����o�7�=�̠�&rI�Gɲ���o�~9������fi�LaE�>_������$|AF�6��(��?4� ��{'͓>��X(E_�׽�Q��Nh�� �`�+^�$T-{�J ���yTU�
�GoT.�������_���/��֏��źT��B��㛮��)�X���!{
9Z�d/ˎ�.�[E,�]��R��"�/U,fX�����-qd=;h2����9R�ȣ{�)Ͽ
�x�zJ����fB#�'V��0"&�0����wr�2��3�2[�j�w(r��^Z�eIK�i��A
����2�ݿ�vM��^�9"��1�V٪e�������7��z��Y�ٶ���5Zo�S>M�s͹��A��;��쳚ob�s�s ��
�O�I�z�����%/x�+/0I�y�J[c_2�f�T�禳j��l:�����yf����<\gb���&g���-�-����W=ܢ���_�U��-d֍��]'��EeE���OZ���r�.���E�53J�1��ښ��ʡ�M��hI�� �D��J� su�$>@�623 %_y��m("��/|}����ɏ|{�u;A�(I���[j��p�l�A��lӼ��(��ۍXvp�ο�JS}p��.R�����{X�aje�Q�O��@�_~a�]\(�+�Z��B�2;pt��v���!�@�iL%�s��p�g\��s��Q:��g:���U������9���"ᵳ����e�g[�ǝ��@�	�/^��(�<����sZʢ�#��{WM�V<����:�����l�D�/���aϊ�*�q�[9)Wil�DX�3{��N����l�QYQY�t�V�V�����h�|�Af/{���JB፲�ˣ��"��^U�׹;�E�]�Sr>}q�G�[��PT'�-!�`��k��.9/;q5�g�>h�OHn�/wv�b��G`���+-�w�REY|�b>:d-"o��Y(��³���^.~�-ŝ`�^P�M
�9�Mr�k�&	���Ӊ,Ÿ�[���7�uPU�e[Rs��q" A��j������?��e���F���RXXEz��4��u$�ǲ�1PV���G"����e}�؆�:����!|ꟼ����w�*#9UU��"�'��qo��g� ����v�w���蠐���֟0��O!4~����)�PQ|�/�xC���e��nF�P���ԁF�B�A�4n�ѦTx�^G��E$�|v��?�BNA���ـ�H��N��^�Di{�ʕ�O��_|�����)�<9�5��Ă�Q\R:"���#?��,��dh���|8�ew8M�����f���x�}���9��_@�94p�'ۥ�j�����{΢�Z��ʁ����Y��ք��:%��^Vk���y�*��DsZD�g>2zj�Ѐ�J��Q�܅�!�����=�a��j���'���N`�l�bj�(�/X�$�K�%R2�B�\���(U�NρUr�f��Ds����Jc�= ��ɳ��b��7|�-o���%aXj2r_�ݭO�CbP��lwO��I��*�1��S>�X+�8�$ԇf2�Q}s�ى��q$;���$�E��-j�.4A&��JYu&�)M>�($D`(~�Z 'WHDw�K��t�;�\����Ɉݵ%ҤLK��x�%�#J����%E=Hx�)�P���7+!�(M��>��uJ�}0�^`��:?O��v&�������1��$Gƞ��u����tH���,�v�Ul8?���y���D�_)�}��!r�o��hJ�'�w��IT��@��h����Lj�r��2V�(e��"D����/w�~ξ=|���mYǷ�?�>w��@�2V��Wӆ���s��>3J.p]�r&U����0��;��ΰio����0c[�԰����nYB߯MK�M��@�"uy9m�o��]�q��r��rإ�a�����K��}^����Ѭڏˁ�*r���Ӥ�7��if��e#�.Z{�?�R�C�S��T�?�M�$E�^�3ܳD��²[�WTndjJ�%@�m��g�R��(�"���-�|e��X��.�	�=�G5�	˯�
Y�J2��8T7���?�� ����TlK�9\�䑴�=q��魛�<�{ ��h=�r���4ύy�Uۂ	��v{�^Jb6�^D�'7y��I1y[ul�~��	ƻZ�@G�d����cw,\��4��.�ksq���yx��5�M`OCC�GŠ�픤�N2��n�q���pC�tЕ>Гz�pl?�4�����bj?�{�,_�|kd�g߿�`��%]�)]hG �9��	&���C+���ك\���/<���V�gҿ��_3���U����m?�m\${�;xKƲ�K7ʿ�o��y��c&���^�fl��~S����{�1m�4�62�C��pکQ�����q��{�s��I�z@��D��Ɗ���&��㥇=f��)
w-������u�
PS
��]�r���[�����XA��è�|��)�6!O�����ٱ���M����l���a�H\�}���Ua&� W�7�h�!�N��^��O��:ad���!:���:����ޝ������8�7 �v�����M1J>j�ۡ��ڒi�s� �3�ޔ�U2�F
���#�5�k*İ}����|�0��8��b �5����b�QZh�����4I#��:DպN�M�7</�q�~3s�����,���p�@1��0s�moz9�Nx�{%�H��3E蓩�_�G����@�kYo5�4\:c&�G˱ ��P\u����ϟ����1���`��˫��!9��"�U�s5����9��ط��+<�w����- ����� Qb.aXg��ܕv[F�E�r��Z�g�E�UBi�ܤf[�8#�q�]����+[ͳ�,t�h7cK�`�\��i��V�ni�O�l�7&�{H f1VpM�a r���x��-o@�Km$R3w}�X�Q�P���ؤf��R�+�x_�R1�����h�?���0��� �����5ʦ;e��WaE*M�+��T�oU�Y8�T�9�D��=ƚ���1����
�n�nx%.���qo��	|��F��9�"�y2��S�T~���ŋ�Yd廨x�lU���G�viG[�I���G�a8��pFx5v顑M,�q� ��O�0S��8�|ao-`�ϢOU�W���C8���m��?�n�&�O��嶖�{�)���^��2[���X�� �1���d���BH��0���ݾј���c��	|�Rcoj-�2UJ2�退 ����5fiU����4́���p�b�:��M����=�
�'���2I�|a�Tw�����)-�z��3C��Ć8Ԉ��-��zoh�tyՖ���[�]�����Co�B<���4R[[�v��y/|qq�Ck����*U��;G��DE��F-�J�Hk�m���IAN�m��\�R쨄
��-��N# x�e�1;6]�[�+��I�\4o�&�]�q���T?�e4��׆����j0*k\�;~�5�XP��}Z;�U�	)���s_�R1!P�V��}��o[�������U�;e��g�4SV�/��읪A�n��7�d�t����o>o����rXP���
��g�6�9JV��Ӝ���+�I�����������{��?]��Y�n�g�$_�N�n�鋺�S����F�A��aLO�ы.�J/�Ғ|�B� �-/�����8	UlNt�G�ȵ��'"9m,�&!/���B�_�7���B{~��V��Q�p����"���JiJ0*��E9,��T��B��Aǹ��X�o�����KE�Y�v�A�����D�8:@��)�f����o�o���C��M�/�J����.�v�RS�ӆ^ ��_�eRA������oj�]J�Yˮ����{�^�]ML]f�4�NUܭ	㝪װ��QWjXZN�D��n'�Z�׉��F�]e���ք���m�-�_�/��o��������$���Z�9�{Fz�G͢]!���k�Nu_+G?. ��V�-_�O)#�;�]4��YQ��ph�o$�JIp������7		���j[J��o�T7L[E2��BD�%I�®;L����S�)H`�vm�A��r�$��K@Gʘ�>�}`�%ީ��qhI���v��mB�,�X݌i
� �uײ����V��*���:f���Py�8_<%�2�q��=��'�?6Ebm�vf �����"3}{R�F2Ȳ��
hO~��v�P]f!����p]��\��ܼo���ɬ����8�G�����X�o���B&J���j�����K�_m^��Bjm�ݺ�jR.�&z���?Se����Ð*#p��Qk�d�w͊x�͈�������TG�o_R����(����3٨�V�H\0l����~}y�	����L �� ���N�k�)W�H�=R�BG��]��HC��}��#�N�+#g��~s&�Cc3G����k��>��KBE��Y�G�|�s�Ը��J+KQA�9R��H0 .��A�F��$Dz�Y=⸡�1g���BU��E����>~�#�����F�rj���o��8<����������E�цi�"	�	�1�)J�_��X�B�]��nh|��=S��Lc`
a�;���W��,�Y_��9���{Cѵ��Jϝ>�}3@�πF=��[����sȃ(R���b;Ʋ��U����l홷��OM�=�T�@ 5U�{���3-��+D	�8�RH�U^�<��@�2)�L?v���ڭg8�w�7B��X���i4t<Ț��2��_�e�w-M�>S�+'���?5
��ٗ�H�˜��Hr�dE�Z�����*�p����}�m�)�q����=֐��W��N���锳Q�S�� ��wV0�rr1�F�Bv>��d�*���@� ��Q��a����.K�P�u]����;�2������w��STOU���P����xy�Ӭ��el�ڄ.���㎐spjxa��9�ml�X�E��I�Cm���-.eD�
�H�=�H���\���GO��BU
�A?l,��5���pt���<��{SY����x4[�t6�[�Śڪv�Ȋ��  �~�G�+@M��׫'�uC6���T���S�ˉ��
����%<���ƞ�$���0�҄Q+3�p3���N���'����/Rp 
5���渾���i��Ab����/Qb=��}�SK��t�8�R��dd���6``�XQ����d �"h~�."?����xU���?x9�a��B>�P�\��kY�:�> &w�"\�"]a��BT�7Vt�
z;{C;��MW��}�����L#K�O� i}uWS��XZ5�<)#�j��Y�-����괨���>Jss�nD�}�QM"��
H�(M^N~�Be�:��^Oz97���%>��>ZU��l�<b	v�_83�p�� �d�!���IK�~�|�Uʝ;���޵]a��zߜ.�yx�>���'"F>�>@��|���C/�fGq�R�U�bfN��T.��`��{�G��_�&��_�f�亟�0����B^�nV��]�;]��8{������r���f����F6$�n��8�*��Օ~ǯʂ��{��xYQkZ���P8�6��W���On�˔�P�r� ��s����{���SP�`�_�����L�J��i���O�C�#��0['��-q���gv�ߐ�;��^e���T2>�S6%���}\fH�,��+RǦs4���~b�w�3!J���E|�,�oElH��L��Z�^�T�~8��r��e�-�ql�֯w��ܫC^W��W��\�S�E?P�D`'}�CJ
�sGN��Q2��L}�#浴��F���{9Ԏ���ޟ:�*6�6��!�������~�:%�k^�w���0dcT��Ge{�a��A�K8��ha��Ύ���T'̳��N�3���|hv`J=0p� 6�~T�8'u��]j�����M���)X��Q�9�&-}�o^[t�����F���ϱ�Rd��D�ݮ��*�E��c��!f���f����v�YFL2\��'��G��&q�aGW�U�>���,
��A��!|�`̿�`�D1���>�
�8�!}L�w�,R6�s6��K^����Ó՜��(��m~�)������p��[��y���=��A��Q{�W�O�8��lK�if[ �Gf�j�l�Ļ#�܅͞��E�5f#�J`��VP��܄b6���twg��A��������t}��}P��% cН��Hw�=��p�nпP��3]�N���j��9�����h�ؤ�(Q��Og��݉M���+����c�;PZ뭧�X�\,�L]��N]�)1��By�H���3�΂�_�s�,�n[z("�4-\��b����k��>!�+
��3���5�J���.ݛgc{SͬP<�~3�Kq�t����oc0��˙ؘ"�	�(x��w�����H+I��O�P���Av���5�X���HY����*"�_,��Z�\��^|�r@{V>)(2�"=��9@���N��^.��~o<������j��/$�������T&�8p謔���W�}	eE���ڝ,�װi���EEN�Wrx xR�z�Q����M�7n���9�9���^�A�[��oV�(k�T�t��6�NwJ�5obȽ԰��e����<Q��E/��`��s�>�%rhf�l��'iD������T��q;�aI�\{�����J�
=2���ǻ�y���?-��<��~ˉ�/bb��JSW��C�7J�ڰ���R�D��L��FO�B��ʡ� �O����4e�I�ݰ!Kv��SbO�'M�X�|T{���*d㎎�|ϴ��^W��{��� ��gM�$`C��Lå��~�&�!���zG2Q����h9Ɓ:J�+Ŗ0�F�BeQ:G�ܽd��^��,�
�B��*��JFK���Y�?�N��bW�ه���2K�׋E�3M.q�hR{ց�x�i׮�.�%%�@�r�GD���x�*�HA��޼{{M������M��w�ĵe�n�m*���^K7���<BU�VY$���Jbzh�g_?��B@�˦{���9Y��s/۶z����3k0���®$c���:X���?З����o�Ǘ3�\����F�}��:�����hGA�ۖ]�ؙrBS5����������6	�4�|��5����� lC�׭ClJ�n����1bt�Ϥl�+9�G�T}���H���Q3z�.�4�������KYt�>5�!����6�s8�|U�Gl��Bq�Oc̞a�F
%?������
�H��ƭ,�h�_1g�$+
�M��4���6��,��@��M�aכ�{�tSH����8�B%)t�dw!Zq���j��_�thH:��2_?���Q��Hg̹���tGY?�ǔ��������BF�۔y��q��!���i�r���=By[������oRŏ�t���,���E�؆��zf�5�/�~]pN�̅��\j�U*�����L!��7���F��F��ǊE8��):ҽ��b������1�.��r�d<��_�,�,0/�5�T���莴P��2�����9	�Ӥ����xc,�i�[}�'w�v�mP�r_\�/��/MH$b��	�n��!?�=5����Ko�&u�Nrq�C?�M�e�Nڒc{Dy ��k5��mz���$�WS�<_�N����**�M!5~� �W<q�C�ge4�Dz���c���rf�A�9ؒ�����A=�?��T�X3BNe$V^&`�b�A2���f�)��K-!�si���E�����]��8�;ǌ]�T��nV�,�%N�^�X�E�wu��]��N�⇳�v�g�g�Q��w2���Q|�V�>���%j|�k0��\m��NX��������W"� u�w�5N�c1')@�}�� ����3�B��u���L�V_)Y�_�I��^��%�~mЂ�Ü�,��2�c�:���:��MX���E�K<��#��h���*�k���§D�:J+�'����lc"��J�x���r�WpL@������j.����7D��w�$�]5d���|^`ݬ���t�:������D^W���	=;�B��{��Ѿ�!�~A�-E,�����[7�m���P֒�;˷ա�&�˝ݲ� 7�NyxۺIx�Hv�(�+�&�W�&�7/�I����L�k�:yuJ�vɵ��ϰ��>]�1\	��k�ۙ�s�I��M��v&�υ�ό�M�+����s/����ދ��0#� M��tş�����OX'��,=]&oP��-y�3*U�v]��	���Υ)��3q�Q��4�K�RGW�ޛ�*V'B�f���r���H������^m�����uඖ������O	z�~�r�c���=�������;P��is<��񛙀�HM�͔4#y7�k�p<��0u��P&i^�"ϵ�"���щ��%��l����v���-�׸�/F���v�s��F�������_�Æ�����{�@I�4AX�F��;����p͕J��;@佤h񓒿��,m�Z/�=?�����9����yݜU�u�u6����vi�"���K���
y}�~�#�[Ⱥ�m���*���H�X�I<,��O�j��o�.�\ja?��l�rLkG�5v������Mb����TOg�o
�m��
�>])��
	��Sd8]���vEvա�~_�$��#9	��B���������Ih�i/n3��h��Xl�6ׇ9
�A��r�y�PZ&}�$���SV��Z�(���Hӂ��k$^ݩ-����g�Q�/ sn�Q(��t�Z�Z���8Y���dh����c|h!�B.Gy��]�o����~�i�4�QXJ-��ӟZ�����ݩs���=�5�N��Hf}�Y�{3hC"���c�f�i�F.*���q7
Z�Ow�|u@�@)�c�wD�Ʋ	r�Jh��<ǴC�'1Gņu��%�z������WI�����'��_�~T"�� ��2�?�j���ϐ� c��u h]`"����ĭ���?���H�]�C�W��rl�	�+k��<��d�h�_�x2�H��t4B1��qM�If���S����h���(�g�uJ����(QKΑ61����+;�D�5���Cݙ|X����v-ձ����j[$m�JԌsU�R�q?cV��A|�e����5��8a�Sҝz*;؁|{��ϸ�K6�V���˙�2�$�Y��p�U����a��Y��h��B����ڿ/V�z�U�^�Y�*���~�[���ly��'F�����(;���o��o����>*|s�Ԏt�Tͥ����cNI�y7� X�˰�]N|��Yf|7��Y9j2P���W����_���U{�8�;�]�����7�o�4й���k??;F�+��5q{sh�R,O{ǀ��jA�Ԓ���fۅ�TX�����P�˗��P��֯zJQ���C���c��&�[1�ģ6|!3�o����3r
�J��d*3>$
��Յ8�ri>��4m$V�e��Y������L��P�` ��ro��^�N�١�)�GG_�v��}��^`B�n;��$��:�v!��򖚙�r/�#�1򢢓�93X�~��"�����Qp��1�(���{��Ý#���7MƸ�g��g�<�uk�gD"6���V�s�*�)����S	�9K��'�����дƱ�"�uZ�rP^���4ۅ]��xT`����(i5��6?CX�Y���#N�?p�}�e�]&�A3䞛Ʉ2��vϔ��d����6����l[�D}��#�Ы��c\0�跂�VN�6�t�5w-�F�t�B��%@��3q�`�A��ᦨ�|e�Ҕ�^�!����u�Y�_}�y9:�|)��Qآ!���s�E�[D��?��ohw��?�X�&0��1�}�5�Ş�2��WO�/7D�YU��I�!������6N����Q�V�=\�}�{��j%x7�j���',��9"�{��흪���@�iJ���0'�����?�w�NH�+!<�d�^�(J2ԁ���5�~)|(�nr���s8�+�)�����*h-HQTu�Ga��V��,���.O#Rw�Ư\GM���D�v�W "��e�'%u>��kc�T{�0�,�GK*��u��[DZҢ�,��ݵ�F@]\������,ŀ�/d��l��K�cG�xh����D�H}FL�J���T m�j��v'�zl�@�K���k�����t���hMQ�-Uz�g�D�)�X�+]Uf[c�dd��<�'	6��&|	�f��ơ�<�_j�쥿�m�'\ i�P�yp, 5wb5�v.K�E����zYw��D��@�A����(�D38CsKHy���5]�+E��h�'f��peë����{�n�+#��Ż:=+�}˸�F�pq#푅+ͥ�s�KE��n!NbQZ����V���@w)���Z�P+ '���7�BkZhR�j��8�"9�cVa���m�;�)E�pt�	�(p�M� ;Y�����,t.H�q�R|��ۄ_>5R%���5Jd�|���C'$:��:��������k{���+T�����!C�gPH
�(�l��^h(|d�W��9ȟ���RQ�,.]�-��ߖ��z2��/�3[�w������!R'p�z� ��o�Rzr��߷ �e�Ƹrm���^mh�x&�]�&.X�����y���d4�fx�m�$��C~�_�#��y��r��mk#���<1;���쨉�����{�X�p�!},?� 9:���9w�\k���9S������
��45���\->�E�Z?f����_��G����*���h��M��[���p_����|�YBg��Pd6+�g���X#�e�s,�y4��UvYԧv<����:�	�CN�KƋܚɦ��\ib�C�bҶ�Q��\�?A5:�hR�7at!������iH!���sUmݞ�L|��|*V%�<h7Z$v��dm��~�ZD���7���gۃ�'[mQ[!Ų�����TXNb����]��&G�@*��,��T7O8χߺ#kLkn�r�'�(ws��p�_m��Ɲ0溯���w��Y�������4.�GT� �Z�A�\mgmN��\]�r�&���-��CK�ĮώB�]�'�߅�!�հ>ORW]ֳ�T��!���qPTN*k�֋>�Ү��_�t��g祊C�_)�{�/�����rǔӕi�����V���ȋ=�n��6��~���Ŗ�M����Y�@�x�ǱVjWL^O���$����)��y���OV=�_Ꙃ�i3����Zu5Z�s��J�ڔSY���O�T�tW��'��
�5��̕|�B�>�N .�Z	�o��>8E�� ���Z��ʷ��D�W\綑ċP� &�|X����V�������m�$�C\��+@f�&ڤ�q���{����hj���V/����%�����U�F=n�S���S����+��=��)^R$��	yFQ�C��nӤ��4NW��L������G򓞣�=�Ư2�e��;�6X���~�̠` eQ���D[��a�/�h?ue��W!w<�NY~<��Dƽy���8���_1��4*��.��k#��\���&�!y�Ζ��T]nQLĢ�N�7��`�'�s|K���h6dC-G'�3ER���S�v��]�Ԓ������v`�5x�q�A�����[:���
�3�2�]��=�Hc2Y�(C�S� �M���-���g��o3m�5	>�`}�{�?;���r���o�O?0�n��켵�d�43��u�a�_����3�<��á�yX�g��%��_w���z���-�w�@�<er���y���"BxC㽘�N`-8�h�\lN��$1�É"OE�A��U�x�����K�eD��T��u}^����b��d�����:P}�4�NV����H��9E���~���ߘK����f�j�Җjɐ�LLء��P�(�"����Q��~�}ƙ�ݴn��J�+vGI�V,<��p�TfZU���v��Y�|Q�RN�tzC.%sXծI7B�����}�����Qg�:��=Ğ*�J�*�O���֝ӣ�I��_���\�i�	y� ��l"=;���M�������Lo�����o��8Ś5��Ϟ���f�O�ۚ��y#���6IV��*nx$"i�zgUc�`��x�!��˫�$�,pҬ�U5���#4戰�	~[A��۰�׵Dz�ȸ�ݹH0_B�{��5��T~�D��鱅#䒆�=���씉�g@�F��B� b(������S�iԑ�t�t�]�S�g�n���{2���e��Vq�ҪG�s4�6#�ދ
C���i�4,Q̉E'�]����i�)v\��~�aW��/���?�/�$�Q�o�|�p��e�7����"xi��o��A��&�&��[�M�{@Z�S�㓺��q ��K�[��C,�g_��P�v�7���k�keN�4m��H����mt���O�!��p���枋Z�B�mu)0����C�:�ȍ�L3�Y�+��:w������"�C^�urX�N�>��
j2O���7�A��+�g��*�/�9}<�e����]�1To�9�4�_ς�&�LŹ�sy*>'�O"��G��AN{�$Pw֦*�Z�~ұ�޺�S�.г�F���垆:��3�*$1\e�z��}�qE���?zz�/�P�o>O��{NU�u�<�=�����f)��Sl���$>�t&p�M�u�FM�/���(A�hNT��L#K�&�ȥ��tG��IM�ɑ&O|6��݋dt�8�;��z>R5�ʗ ��-�Ԭ�J�:O?7�gM}°��Y�\�~=�3��	~�r=wjt�3��y�J�:��%��B�Z�Q���?T�^z$�����J�0�*�I�g�^7��2�:<f��3�*|`���b���hH�S̓}7r�(�n!��I��j���*:�ڙ+RVvv�	:���R�z�ө��&���>� ��JOvU�IX�E96��:п5r��[y�8z%��t�����d��-N�B��]�I.�z2�:9'^Ʌo8C��V��M=�J)���N{/`�(Kn�:1`�J��-�;g$&���P>���Y��΋uf�4�5���U�7�ګ��lw�6N�+(�G[��	�\FZ,�qlľt��?��C٢�J�S�^�4����|ʻ�w�%I�"o�(���+���!�bв����u׌���=�$����Ӻ��p��ZwF��c�gh�BNJ�0ߧo� �9���mU��`9��5u�9^V�s
�dI��r(�3����uu���R�FM!Nh���o[�n`�g�� ��ݰaW�IY���y���v�۟���}���`�{+=� �\9Ҍ��R�s}�-��w���^w>�u�_'��|{�+PGZ__^qCe �d�\cmzg�Ŵء�(�s�Z`��ȓW�۫6ķ��w'���S�ޢB~,�*1Q�e@=d�P����?>����Ƹ���֓�O4zDZ7&��p�9Ψi��E������p�n���O����O�F*�;y�����o�o��\�Dzl�R[�{������&�������Yy��8^��w�ϵ4.�2ꇦ��F�gq��}��:pz�a�2[�v�|7�iIF�Y������O<�"
����(D��,f� ��1��kQ3FU&;QS0��\;f��e���V;J�����ߘ9m��&��z|�|a�}�F�M;�l�a_�-�\E?↮#@3�'}L��G'o�8�,��]������
7��4G�ژ_5k/���"����ҷfvӮ(�!O�z|
�؄�"���]u�=��$��g�-�Lxz=���DE�JAU[�b�I��۴D�R��\h�Ҙ���;�6a��,�`�gwb�7Cs骴��_�|�^hAɇ���f�o$/V�a��YB�pB����D�寓��س �"���,�59�Χ�'_��eM�l��讘߻{&d��G�6�fe��<�5g|��N�Ԕ��O��2˖
y�s���A�WK���d9��H�+ʘxT��RW�	q�3�|���w��*Ķ�5?�AdZ�w����S��E5I!�0�4s.�s3'o�k����B�(����\��+ht��,�y-x�(IL&�e��z8\�\� u�|
M���5�Dۃ�E#zF ́W�Z��[�u�^�����\�h�sEd�C����H�����J(h9I�'�_�+'�//E8
̷�#�G�#�?�s���͹�U���\�8Z�#})���E��H�C��\}�n��e��@̽J�(9ȳJ�ԺԎLr�Z�a�D�vN�N\s�L��4z0�r*�W�܈\�"m5Q�t*T�Z�3^��8炰~����Mw�{�1�.n�k�/D���V��&�&]���W�Ѥup���ӝ��}���l��<����/6�ڐ' �s�7�H�}�^��N�=Wv��KK�����;[�5:Mk�}ĳs��������w)��<����U���PRiX=�b���6�p�8c"���L�-���1"m�N�T����:J���%1��4✌G��>¾9|dj�rx?=����l�H|J�l�P�"TfI���zγf	'�F�[�/�����bݢ�i�@h��:XZN�F���=�����
��1���pw;�fS:ҢNf�XT5EpP\|�*\��wYU���Uf|XB���w���r5���Q=Ǵ5���Ӷ�4*���h�p�Jv���+S�Sɞ��s hՂ	`��d�.9hVf2����x��1g_3B���W�V�\��*����-�?y'�N���I;k���O�;'a-�fW"���(|���Z.���(�O	(��s\�O4j�񔑪?;m��s���T�Xc��ߧx��o��u#�<����l����[�������Y�k�煑q��;�N��\M;�k}��R�o��C�qz�y�kO�1,pee:��}<���Kͨ��D~�����GC����q�ҹq�Z~����xM���y�*��KR�.m��(-S����£��-8A��'�
�1T�S��Ϯ�SC����L�k�Q���D�Z=��pڸ�������e��&(���5�>��Y���ypc8�kʿ�?�eǓJ�� ��.:M[Iu�羽�Q��3`��?�~�2����^�F��,�\�Ԥ�!g�\Y���{�W���?E{�*P�_��!E�:6�����i�Q��wȬ�o���6���"��I����[\6�}��/H����SA$<�L7�ȟ7JLk@\��asj���z��y-�OcD��l%ڠ�D�ߺ�,F������V�sݝ���6� �wlQ���q)s ���˰�5����`�׆���l�Qs+���"����0"|��B��zgw����	�,"��!2�`]U[�J�X�|�<��ȱc'nP4:��)���.ƚ���*B>�[G:��?&�Ñ��{��v��U-��*ڪ�Kh��]�U��V�س��j���jU��P{%v��=b%jDl����~~� O�{�y����h��[=�zo�4��D������b�O2�NbuŞ�)�9������t��e��\U0��h�⨒	��3���{�Л�����ks �6hS=���*�v?��{�kjaCg��-�f�H_ST>�����w�qD��5p�uA��`Eǵ���dkwt0��g��{�׸!��YE-�Gȷ�R��4ݩ��௅Ó�,�9�S�|S��h�֤Dc4@>�*62;76�3�עy]g7��n�,[ߏ������1X1l��MMA������~��4|�ƞ1`��Ƌ����^b����>[�6�cM|��z~��c	�0)r#���}�����[���m:w�`����}	�*vI���H�*�W�J���P	���B�E�a�gK��f�p9��xJ;3C8Sq���?~�~�8��ąs���+���՛���k�kK-��rr*Ëa��|Ά$<喪e�o��/M�O�q�Ǿ�Ѝfn��|fW�[�f��yϨ�bʈ:��Mz�1��-��z;�·�����lr��4�x	��y��%�[RpB��Ew�7`�=�Y�GT�Q�Oͪ?&
3���q)|ᵣM]c͓9�� ��T�&�f���V�0�R�x����X�-,:���&�ʤ����Y6���G�Yŀ?�YD��&d��}�q͝����n�2�0������<d�����U?Z�e����I��#��̦�`Z�8�`�1��1��d��.�
#���_��9��6*0r�JV ؈��(H���ɟ�����:�eS>�l*̘hQ	�Z�������7�;F��I����W����sn���
=�����6i�9z%��_��h��}hpG�3�� �!�� K��`R<�
����F�4�b����(5�W�I�\_Vw ����]�{�+��Ĥd3'ú:��nnt�-ʺe?83i/EF��}F)^\J�ס��[�Zt��[�*��#�0&x��m`�d<rū���| `v�Ǭ��qhs��4H�x����g�#���=�O��1g�h����v�ă����Tk�p)�׀��j����e}8��,^O�I~8�f�<�X�m��i����H� n����U�������S�����{�[1��Q�xU� _`�6�o�Wts��b@N8�j�b�R�B"�ٔ�*�s�<-�%�:����n@L�^DGr��_L�	4Zȩ/�E!���7�TLd���gtq m���Ƕ+�$�-R��f�Ӈ֨�>�z=��C#8:�%�N�I���� ;�^8�J�&--4{aZ�����W�d���N�Z���K޺4��l�;|�Y�af�W����
;f-*�d���۫R�y�Ç��-�4@��)	ZI:e�]�2X���S�{�Q�����z-��:�Qܢ;g^����vU�p\�#r\�9+�3!����������s.����[�Rv�-��JxJ�6����%�'V�y	n��F������[av��)��3��%?��֯\��=�Y�J�4Q>��_/��,U��z��̀��W ��T�����\brK������	޴��}��KG\L�@3��K`�X��rxQ���3��ϼ۾��&�zdhK��U1��V9+�ՔK��BN�!�#bh�Mc9:�pQ�?ֹX1M؛���{�a3G����S��PT�O���l��w��W߲��;򽏹t�:ud�5)��{2R	�v}@�z���G���v/m����bQ��e�"�q1��qQ�W�7i�1Ro�C��ʐ�!W�4�Z[;�6��cV��۽;[{2�I���=��)Q�9R��̺��Ӛ�R���t|�,�ᇡЅ� �B��V;��a �+pj4�B*�}��Q�!�$DM1�Xeq������'�,���φ$7�9��e�ΐ�k�M]��+e@����ȴ8g��~_#k�Q����>�k�Q�k-��"�*�s��h������Xf���'��r��3�
�	K�rb�T/KJ��������E�MGp[���X%n�γms�Xb�=�'��+���3�A-��I�����l��"8��RY��,�i�����e�,�%�����N�=aP�1lHW�i���k|��p�I�eͱ^���:h�����Bq���̉h/R�w
�7��I9jl��x/[?X�S4S�㰃���n��??�� �j9�K}���<�`&�ʳ���6����K2�-:)?S�"	cG�+�U��%t��G4A���G� ���"ǚ�H3�_B��ӉH���g\����=���؀��[w�Cuts0dgok��|���(����8����F����7��2�fqT�A�K2;�<#xs��k�?�TIS�ݽ��a̹\���9��lѫ�88ON|����&��SD�k��+�U��yS|�����¾�� � �'͒�,�`���5�Ԯ
�]�BA)9� �R���RĨP"�:/3P�c~�j�i6����M\����=P�ΣY���/������S�}#Q�}?i)��J6kyן�˛g��o�L�s8�_#�
�af�ɵ������-� M�L٥*��W~]jB%��J���~3=!Z��
�q���"`ڡW#Z�]*w���mYuO�� �{v�����΢q�sZV]]�g�޺�wa�l��9J��l�ٚ)��T���,"a� ^�E�2[�9Q�,=�� ����w�X�g�8��m:��:��b��"�c"����[Zb��HAK���=Tw�Y�q*���R�- Duq��!�xR�����y�z�93�n����ҹ�^�����iE4�!���?�^����V�s_��J���E�cG�j��'����
I�JBAV�k3̓�/S����K);��~���n�Qe����� ������/YW�Ŋ��=����&1IHV����BCkk~p��}4�!�P�}�,e���¢%�����O7s��.�jx,�<�n��J�c@CT�4��l��~��UJ���p���'�n+�̻�����Y͑�r��� ��4A�'��U���-@}̲gk6�>�2�BK�,�"����	4���ъY�[��%\}ɚ�j��S����Tuj���Ã�c,�-k�[���2}W�7�-SӃ�&��i.�����ImL\P<�9��ͪ��K#�J��z���{O屛M���1hs�{%����-�r��^Y�E�QI1�$���qE,u�	^���4V��ތ���הt�=Kڱ��%�&��w����] z�����9#p��ί1HJ��t��jF�n��U�����$gs%iWW���c�>�F#�l�-�i����*���$��0�z�/�>�!����M>��<?��]/M���F|� ��?~�᧞�����j���_��%�����8Am�{i�3d|%�6yWn�4�$�$-�+���>�2�/q���Q�w��5�cMK�[�Q._f[y�Ks�΃��q6�M�ڂ	6f곘it9Oe���D/|��3�/O$V2l�=�O�@5��ns��$5.(j���N3+����C*����>���5+��yv�_��)J��I���S�}���x���'�T.�,���R�����z�f�_��u.��|F0e�&��0|�~�f�O��
�T��k�BeG*2#�N�����Q����m����h���?���y^(�S�?t�"�9d]��~y��鴙D|�}���UޥH��S��RA¹����1e: 8�&��`�B��5��GZ>�U�2�����8$av��6�р/��y�%�6�\c`/��>'4�ܹU�6�ڮ`+کhּ��Ɖ������bFc21���RD�3�0�&HDD"�3�@�?V� L�'�oP���$�qTolܭ�V%��tq�P���V�g?t2¥;i� "|��8�z�㚺�U60[I��V[�
�BV������5�.5����/���]�>BW�*������x?q��Mbp����8���\ciV|����[�-V�tFKC{���_|� ��j����Jϼ�1����g���w�W!F�d�qL�@T |bQ\0yog�r+��^-䛝_����3[7�e�%O¼68U��W,�����]Q^��B�<��Ʀ�p~���H�3�њ�u��L��+<)<�X}PT�$�UY�f�x�:t:)�"�C�"�ޡ�E�~�/D��/Y�L\�Y��0��Y����f��ҁ�.�ܳ}F̂s�45~���뢒R��1.��'{�{@\#4����P�{���}Ǧ���C.����
O+E'U�m���[1��I�	����gh���TPE��;_�c��%�B�Ù�p庯�����ގ�.�a���eS��L�P`�,+O}'=���@�Gwi���)�Z�l%.-e%���W��U[k�8d�Υ�.�f����T�kರ�Ӧ��!�[[���D�����mﯬ=fFnmcX��D*N<�����p�LDw%eIS�Zt,��_Eu�I9x�L�pF1Q��������U��k�+��Φ����Ib1���C@KT뇓=����q(�Zv ��k�u�����L�>n�s�KP�:��n%�[X��l.m%����q`��ӽ��»�N���2S��k��-:����K�V��j��Ae��B{���ķ~Љw.R[��*&\e���� ࿮�g?,�m,?�h����U{�,\��5=7�3O���Ml�y�ZVV��bo�Z=�e|S�� cג��?D��V~�I��J/h�C�����v�f-���m���ɏ�R�q�睁J<(�e!U�x)���f�)U�g��(]�������c��pO�cXRg�����Y��2�,>�f5��K������M�`ݵ�_�R�;I�m�7֬�WQ9~Q��w�"�$9`�����
�lB?W�H��v}��v�����h�>l�X��+�-�REE� qp=4��+04I{|R��@����&wﹷ�+���r�$�g�R�8�o�n��,��t�!W��
ٳ])x.�k&�\PuZ�8Tr�,�[��͝>�j�#�<u�'�л�d8��ф�b�4[_���p�ީ�_�h[&Z�]4m��k2@u�0�_O����}w��:ȺC
vK��ʺ� ��"EwNA�`��G`��-�V5��_Ńڟ�L$h:<�? L����Õz�+����cS�RP�-2�y��WP��1�P�;ٿ�:�󘍽 ����Us�~��ma���E=��>�B��I�����u)C
?\�´3�{�[���.�L}G����l?��f�;��%�h�r�%9��sm���m��&�ծ��n��"1�B
�+��pT�t������W�h�z�l�<���Y���ڪr�(�W ��T7d�9�	lM.�Y	���R" VHJJ�Qwo:�d�M콅��P��
��l��? V�+��ț=O"��l���$�(�Տkyߩ�#��3N!�1.��r߻Q�� �Z�7Fny�t��`����R�_�:-��Q_���x�Xg
d6�<�e�%m� ��M��rN��G:_QPOW ���DN�x�(k.��DwC��sQA�ӏns ��U�0]�"��������Lώ.)�5m��F���Vm�T��W�I�&X��:z);:����BT63���.���������-ɾ���az��h�v&^�I�r{�3�`x�|�E#��e�+�s`\��|F��ʄ�gaֆ����]F?��X���Y�i*�!x����H���S���֎�����7�`!E�-�u��dwM��=E��~�N�#�i��e�$�s���,��D �Kz����Wk�by��_TK6��;F{dg��b���J��X%�Yg��x��{%�'���@6f�w�� �w��	���$�g���+ �
�A;�K�8/�<�2F���W���&��@<_�xl�(m�$�[(컖�]!���u��ص�Ë/ī�ؾ�OZFB���|,�s4+f6�~��Od^(�Y���P�ͻU��E�jb�GÚ2�Ng�+����-�W�0�c�^���&ⷕ3	��	��t���T�M.�H�6s$���c�F��@V;w�3�)��^?i��Mn!wE�w)��Yu�r�'�48�39p52���W��r��O'�tU��f?:���"'�'5�T�	�їk��8�J)�4t񈔑7������R1�%�y[|�]��Uυ�1.iE�RDҷ��9�L0�2��ro���}qy��N�'�c�_��y�K��T�1N��g�g~�����)����z�m��JyZU),l���8:���J��fb[����(�uS'b���ԴF�{Dm:�9	�C���n���67��A�+8�HT�r��8܌ѐ��,�:t�/,���0�W�����;���.�q��<�{��1�5��C4�1O�.2��9���I�z�o��<��3
e�rc��QE͒�،�R]��j}S�k���Ո�c\�\��r���W��P�y��'xEZj!�vLQ/J�1�����tSBh�"��dΚ��!|��X�܊)O���0�'��}σ�Ӆ1���{���񼪔�S���n3���5��R�ʔ�����p>���z����H�xq���.I/��Q�<b���|�̬{���xi�q:��2��;!w��UޛּN�����.���]6�����Ԋ��_꯴�{�� _W���c#�@[���C�D���"�����:-J ��c�I���7E���J���P\^�S���Tc,�0��š��㰴9�(k��X���@�EI�Zp��O�uc�(�<k��}� �)>������TLν�Լ/�
lMi�q��<΅~���~vN�}�:%��8t��ߓ��������.:��Sط㶔ge�@u�B����)����1f������2�ǆ�e���kq�_��v�5�ܼ͗�ƀ�"�Y��?^� n�m�c�������R���o��] r^�˨Da�g�E�^`@Rjrjo��J2�0�J�o`/���C����y�h�ߢ�)�J|��:��鿋ۮ�
<K�ͳb8Q���]X���.��Y��'f�e��W�NE���|L}�RI��M�s���0}1P7{wg�/����'���O 2�WR�:ݸ+���u^M?�x�<_7ܭ�s��2[����*�������6!���8���W�!	�f�g@���u��lw���uo��i�&�l?~
�[�pB%2�I�8iyt��=�@^dVl�����$J0��%�')�ʋ�܌�8#�������S X�N�����ιa{���}&Di���i��	�7_�샥�9�������zl]�F7�p<�Ì ��g�h�/���s1w���Ǯ�|��4GЊS�l�`��S��?K��z�2���V|�^�h�ï�+�3�5��wG�8�M��>��{�o�{+}��͝��K��I�1�	깫��9j9@�?dy���"�c�u���*Pj��v8��[Q�=��1�r�²ePAQ��m];h_ykP��E	�����pt^���Y��ɩC\8xO���Q.㧫�+q�t�Z*���df���0:�)�[� D�T&*���9��M^<4���ś�����[�d9HNC�%J����$l��p�s�W��7G!c�=Y&@T�wr\��̉�s$("P� 3)���D%d7 &���.}/%R<�h49������@{�ƚ?�/�^v,.� V�ȦQ���Z�i6?-q``���ڋ�af|m����^'���'�M�]aXa�� �T�Y�m�b�kF���µY���N�TО=κjRa��
��P��U�p���ǏXߚ����U-�C�ƓuGs΄��]?Z�s��W����r�Ow�
�a�����?��M��%����@9�~�e	Eij� ^��\�c���_��m��N^�;u��S��m2B>��M�##����Z;i,���#z�CIq��o�|��0o-�L�@V�h��&����_5:(����������kq*�E�'��#U`T]Z~2}7>]�����&��cK�=gdH¯r��^	�%�h�ŻsR�s�W�b&/f��;�$�gm�<��O+,{��\d����㝒/�C�,���Sn��IWU��$f������W�ݿY4���ҾU�HBT O5߫�r3rs;`�R���Κ��вF��4�+����u���-r����ť���=��J����ogI��;M��VET��`��Y�V����9 z9�O�;���v藑E�ԺiҐ��4ϿN�.~
ҎDp]`�p����&@��Y8Рj6�!�uް���L���:�ʝiV��A���S��F]^'a$����!*bY��|��
��R��J�8y������'MSsM"sY�TK'�=E&���c��������R��ܽ�6��3�4��LD��z��y�o�<]��S�X��$.Tt�VI���6wI�z����BG��J�-��F�'��[����>���l�����X=��L��;�����q6+��.k��7�#?m4����U6��1�O�ym�_�,/�|�������e��C�0F�P����]����|��s�����^�K@�J:�`�3^�q�
^�6#��⇣M�����m���H��c�č����1�&7~И��2���ԯẄ��t�8���M|��W��֊����%^~�ط�Ǎ�@����,|�EL�K��M-NE]��o��I"�*v�+Y#[��f�y9es�.�^�.�h�R�\����rr�p�������-������V=>��rH�=БƊ�=:ݜ9�?�׶ω�����_�BZ>x}��p�X�)��B��N��R�e�B�H��<kS;�Pd�T�H�8y�蔈��������wؕ��J�@V���zED[6F�(�[�b&�V�N�1]A�����e`�t����;T}�\]4�o�%d�g���.u��3{��mK�9��@g��m�Y �$��:?t� ����ú�>�CER�C��?�����P:�#Y���k�C��簚[5���n��-p�:�9���NQh =�E�ͫ	-��>���A�,�}�(D���d�FM�%^�����t|�'��]�*'EKrf�g�L�܀ҩ�;�k
�k>J-R0�4/!=�Ey��Ni�	�n�鮭�@;��s�sY�NO�)ڮѮ:����ʴ�2��I�.J2����`Ӧ�֠�{�""��EV����w�b�9�Z���	y�Z�>����;��d��d��M�Ѵ�&{m˦�MEI��`��)Zи~�xI�
�b}�;���O �i�0ֵe�|~��qv�'�J���7�}քsN��+mcΥ�RNo������ʪ���P�����2-6L�G��[
�W(oy,b�N|n�kF&7�������j��O���t�?�E,�����ʙY�;�hB�|$I�f�iU��|�:F@,�����]��쌜S>��l�O�]�y���?�t��3^��pws9[��n]1n��J�o�|������9P�!������G�"�Ȝ)O;G=������떴�	� k���O�.W1�����l����i3�u7u�\�K�p�W;E?�Ă=��T���^�z6�(/'o9�?Ԙ"s&T_̼Bk/�<1ra8��9�5 d+	G�	�p�����B��lZz��Kf�o��)�P�� �����~���{5�!�
SN���a�k��[����{z#ZoU�,�\|�«t����Kmr�U~��ې1^%.i��'5��38@���.%9N$+�`�{�p�i+̈́��P�rD���Ӌ�+��
�����M�HB����c	a�k@5�e?�%CȢ��L���`j5'���v��8����e]j�N���+��r ��Tʞ,�����`�q���|j�-��@A�'�[=o%.%��?�K�p�ZY@[[��C�Β�B81���礩>1�����ƨ"�~C�T�p3rk{�����f0>�G�Tйp9Fԑb}�&`/��oB��oC�$H.�V�p���pZM]���#YOH�A�0����$��1�͡��_mk�n�'#�SVV�_���p�8�_"ڢ	j���a������1q�84fLb�(TO؟��ο��t��݈���P�g�|z�YP��[�&�$��nq|��+>r��D�����q����
�%aGK�Ec:�/!j���1��F�����!�I��I8D�K�Vg��I�a׶�2��\��:/�2m�9E��Q�y�zu:��� ;�qOW�K�J���p!ݔ�hϵs��ɪQNuw��no����îi��1�d
D�a�草��5�aGKb���`�]*���Ѕg�������*�rA՟�O64�� �NІ?!��|�+�Z��OO[�U��ٵY�X
-�{��hE/�L��Ǌ���=s2��}������7��jF��	ڷ=Zc�Q����|�@Br�ΑK؊����>���G�Ȫ��X�{c�~ ?��7�!��Eq��݂��L�F�v�}���|%�y�T��\<n��
m6M����ur�b�g�?�cQ�D�+;\���L�|�K�]�Y��x.�1�?��A� N���n��Oov������I��#�B��n-2�*���p��~o�Q^���0m.>�
Z_(jf����*��d3��1��5on��K4����Wܽ��+@�4+D��٪��0JKY	9���:b�źN ���\����:�9Cј���R���vr`�ׁ����L���)��i*\W��G܇����v
�i��疚*엠Y�`�,����w�E���ѐI#�;�k��:�=NP�x�?Ґ�g.Fkn��f^X	F.�>���={S�4"o�'���Mݷ�(A�[g�R1�|_��q�"^��^0#�xI�[�����嚸�9�3g*���L�b���S*!8'�O���%��>��ȭ�T�����j��@4�W�#�'���x�O�f������P�5�BϊF8�ok�Ļ�2L�b�f���� ��D7�����A��e�9?1����y!�Lx`C�é�î�����1����Յ����e�y���X�[�%�[�ϕ*y,�=P.�{ ���_��u����5���tm�g���s����,�B�3h\�w4�1��H�����6k���"��%��g�#��.jx�(���=���3���\<zPT�����e<7�qs ���ԡ�O��_2Yd�WN��9�vNG%�]�X��'��&�J���-�I�;�O����]!��
��y��WAI��Z�Ǘ(�~�g��F��B�=	U����^p��|\k�s��Њ��(E!^��#���m�<�)�?��?��;.�{��d_Ӱ�쓇[9t'�;z��A���&%��.\���(�b?od����/H�t������#�w�wf�@N.oOq0+���̧��E�iOw�ix|���Iv��t���Mty����Q����^EܭD��3��}l�1A���nԭ�J�1�����9Z���/��x���g�js�k;f�p$��ׁ�u�U����q��F�-���MKO��Ωh{ͼ��n.8�dDZ(���˩�����G�b _��C�hڳ���=K��1����V��p%D�B��
yEaS�5���Yܰ��V��>x�؜#A��	l�9<��E�c'ɲE���� >@����|��F�l�Xb}T�$�'��:�u�'����s�#X�����Ԯ|4��I��{O��h��V�p����@���������q�An�ȼ�g�^�m�b��q��Qsj�`*�����E׆�L�31+��}6	X��
�}�n�Mi�e�,]
����NH��.��Ԣ3��J��s֟9_�`U���5�kv��/��ԁ*#�R��]L{mTy��<���#��y�z������"��$��mœ�������.������'����4�E�}�M#g,������=�$�k=UVe��y\�N_����eMsU���[j�`��,��	'+��D����&G\Kϩ���q^��m�LUM?�Uب_�ⷽ�"����Л�+b�`v�򩂵���Ww\�ۨo�����;װ5��Q<>�/?�N�uM��RY�/Ն�<��p9���tl�6��Z֌N��']����|߽&g��kj���=\-P2;u�B�AJ�Q��7�m앥��,��7�Eʂ�C��I�i*�6q���z�(�`kHBw\g��S�c�Ha��P��7���wv�ˉ9��ƝwJ&�V��w����Ѷ�Ǐ׭k�����Y� 3�~�k���+Mƒ±�/q���s���?���a�?ޟF,˃	ϯ��6�@��a��՜�-�a���6='qf�x~�;�"���]'#Q�4c|ћ�"��m�Ґ��:b�s���|�_�Щֆ7*I��N�^��nt�~Vv���G���r�Ȥ.J�C��V����J�C8�K��'b#���6@t��/+Hys���3C�L��4�T�>RA��$f �{sqY�F��o�LL]�����ׅ�N��Y&�;s�mB��cI���#�D� O�$0��fl)I[K���o<Y��l���m�6���'+�g��z_�Cy���ڔ=#n��Ǚy�%	�c�[��n��O��	��|�����>޶|.N���Oҿ�s_�~��J7PUUg�H`Ѯ�F���3�e����W��'�<���r��a���ߋ�^�#�!��Y	�(OS���*�F��s��K��9�ml@�����bx�I5�&�	~������HpCʯ���"�Z粤�H�&^y�l{x��J�ڍ�v���^�� �3��o�SĬ
r�_�p-�������>�Qe����Ƞ�?�ou&)^�ѩ�[xӊ����z��1j�H&���쾫�V�<)Ev����[�%5	Ϲ���~xd&�B���l��ڠL2)*��;)8f6�CӪ�}��&ȟ����$ҭ�X%��/����)�|d�F`��j!�m��k��md
�K��l���_3�X�����fY���J�?��oq~�⯧���3%�����(I��lq#$����ƕpHEed��ݰ}�Lmj�1:�)�&,ܧ޶W�2=��ER8J\;��L�U�������-�Y`4n���⓵ ��@����N�e⏊A�DR�	�J���dI�n�����-��s�}�*[�(o(�^����]��#�KQ�;هx���Á,��D��Ot���7��>WW�-�SE�L}���|�dv,=��������>Yf�λߓz.F���/��-�'�({�}���,��́�~��}�:�*�H.�-�Ӧ��N��~�R-��?c�Xw�c� i}�A�U)�9W�)����5�t��[-�Tc����������u�~v�����X#�D�^�f�gŭ��1Ԃ�h2[��i�hA�Y�G�������=���SOp��柚��μ��̌�8s��� /�ORd���*����݇��|x�$���pA��BS�������+�rD��D���Ki��&�k3gh.�s��A)- q�� G��Bq?�!�ǽǿ�m@ܴ�L^��֖�i]�ϑl[_-丌�_�̏N(�rg��"�J�4�-
ʆ?m����q
cl��F\���_�ߤU��M;S�	cG�	�k2��ٕ\��|���mv�����#_�E����A��5�b��-X��qu!�A�G���>���9Ţ%c32�,�.�S_�Z/��ћ�R�SW{l;'��{|>'F�pC��O��Ry8�/T�d�ߍ�\����ʄ�"D�L�G�9��`�9J���y�Ɲ/m�}�ݙ�e/�o)J�\Yg��}~.��!kZW�Ka]F"�;���bg���%'��Uv���On��z�m�;�PmC-*�����A��A�A��V�0�wK{�z+yJ���ҧy�̩ؕ�������L�D#r8�?�S�^f�`N�*�'jn!+bK�v+�� �K ��Ǖηg�.Q�6yw��G9`*�kԼ�8��ѭ�юz�����q�\Y]d��a��bܘ!y����sj��K��͛:Ʃ��6�nH`������;����{�0����n%�~�R�^n#�P'��z'E9v����c���n��`e���/��������}R��B4v�;=�D��?�Q;�]�
*DC�F��g�ݧ��o;� �:O���,>��*����k-/�,|E8,��f����+�v��-#�`�!w|�y���MI6O�n��i[�q����	oA͝`R4���k`&�p~��$��'ý�"�5��ճl��v>��(�<�D����}�a��O&gw5N��҃&�#}�J{e�~�� �>uOu��QsJ�8p#�]�`ݿ��w�xԟ]�#ͯ�n�Z�`W��B���y���/R6����8^�-_�)���`�/��%!��9Mǝ-�Ď����,=z9
��a���'}k���'hC�ס=a�)BfIc���_c��;~�͏�1���m�ߡ����d��C�j�y�R2+s��Cr�����AnYt�`[M\�sUz�vl�tg���Bn���D��˦�,K_V�o33��]aX���2����=r*,�����f��D���F}���B�G3�0��k�.�����U���]�N�C���7��2�н�Ý���|�kw���V��|��^�k�l�جf�%S��k���P���V�qg .�Ǒ�a�^_�W����=,ϐ���Z<˗m_J�kE���Zp���4�B�q��q����<��ۜ��W�+���� �^���"d��$�͵�K�i��ʼR�BH�S�p�S��l�z��0�͙��M��]Nd"��ֈ֝ޗ���+��;;�?�٬��۲��Bx���m�ɝ��� �W��f���w����:x���Ƃ����3q���F��Ȯ��h��ac���Ӏ�fgA���Х�.�^��`=��hH��}�Io9���<,U�0^��m����Zw�H��֦Fi)�:��=A�>�ܛMO�&_�����Γ����W/z֛n T�waE��:7���
��)�������������8#�>w�$�d�o�&����ؑo#�A$("�uP/�����`���s�	x�3��~�E�'ݾ-ݻ=߳�X�XZ����[��8	P�ֻ�G�u����f���WL�`|ɡ�ey`*�e�f���`�}Lf�Pb��7T�j�b�3I �gn�Vh	��Ɍ�S��fH5������*�}����/�uu~J�_ͺV���
����[�����;@8A�jQ����L��^m������&��L��	� ��U��{SG�G+0w�{�J4{��W0���k �rZSd�vF�,��9xN��
-��=j�d�w��lw���U $���:�R"e��q��wʝs�Ό#j��R��,�λ��a'�����>s���[���zi&�����|�?�k�"�c���f�w���q*-Ski��H�@�l�^�?���4�~�w��{C �@�\� ��83�v�.�mrƝ��C�b�5ͭ��rv?����T˓�{����,]�4��S�����ZO_~K�L��ڳ�n���ՀDR�{��[VE�x\�>"#��~�uq ��N����ovf����*�L�v^���ƙ�`&`�����H�?�� �o�*��i����JӞ�JQ1L�%�t�b�|ՠ����q���\�O�Dۿ��0����.\�� �>6������EFb�������-U7���bXґ��G���[�Dlxs��T��&sgv�|�P߶�G�=�6�������&g�,_��|�L�����}���+��iT��VN��x>CO���D��ew&[�J]G�������Aɾu;�Պ;��6/�nZ;](��|$UE�L��',�#I`SÁj3ek)&��Ɨ�o�y����+{�O�(S���gl��s�[�]I�@ӷDw�鋀�6h0�<�Փ��O\�������d���RQ�
�2]�@Y2����,t���"�|�cKY������-�7�������Y篖͌��X�q���4.�&Qs�q[xB15�*�p<�[����^�;�.�����m�Qnr��^S���������,{���Ԟ�QDJ4�c��{T�r����Ʈ�vbt�㏮@����Z:�-���כt�����~F|�4�V4{++�X�U�k�8ȱ�v�.o5n��Ĕo��]���;�̯�L(�/]��ig������T����k�Xӵ3ϭZ�;����uG��@%?��wD�����.P�rw*��A�ݿ=�(O��hfK�F�7�r����
J*�t%�8p� ��֫NߐD�C���s����Q=/��2���P`2d�prA�":�L�*���
S��z�d����nG��2;�T
R��E��#��eOOh+��H��ܜ�a�^6�	�;:p�>�E�[:c���$l�dr����:�����:�0?{ˬWZ��ǀ��IJu�e
�䤛,J��Nh�D��?��DY	�q���]�>���nt�92�\��p���{0IRn+�'���m��M�tO�DWe��c�;�^��o�mu)Zj�R{T)U����lkϨQ#$Fc�h�j�[���AJ[�P��H�T�������>���s���:�9�ysԽ0"ʋ��p�rʹ�{�=j��'w�;Ü�W�c�~������5dn��S�4z@(٠�m�o���ң~�7F�^I���]l=��:_5�1�S�j��4��@���8��a���]��CA��eLN���x���$�}�y�Q�����WˣJ�V)�R���n�o_�pgK�{l�.:e��bgX{�b�	��<2����m�񬵟�T�\��*�'��aG#]<�d��G##�^�_]�{��-2�;?�q����*Qk}q8#$��-�f���D��߅�3�H/]����ڠ!���m���	��yY����$5�XƄ�!H���Q���)�ClC�k��'�L݂l�$���A8a5-j���K�L�N	�|i���d��R�Z^i�d����J��2A�����[�y�`��s-�H�4��� ��i;��$3F1���Lߋ��ŕ��z��Ɋnw��4R: �Q�L��6Ќ��z��GA�G�n���V����ب���y��Hn�oMlmWisR�������U����q`�5�-�����`#"�F?f�u�*��va��s�%���.W�dޒ��*���P����U����Ӿ�L�1�m,;�#��B��������ooI�����^��e})ч��1)% GU���&|k� >�~� Z�,�erZ�Ua]��[PQ�UQ�%zď��LJ��:QNo��̥��9T��gϚu<�y��p�S�Y���4�I-�є5�ϣ���B�7d���X#��&����������y�iI�yW.�#],`¤�^�C�����d��)��>#�6=rٸ��c؃Dߕ�ǑN�.ˉ9V�n!�blq�{r�2WA�ȭ<�:"$���vg�W����ؖ�*���ɣg�� ؏�"���4c�D�cm1�Ƙ�d�|��i�T�|��ҙ�"��n횢����lߝ�p><�Q���s`|����*H+�r�����v�ֺ㷳�k^�*�!�C�����0�WȻ���M#+#B�'��:���E�#���l����Dt� &/Xҳ��ۿ��y��ICJj�2|����D����E���4��1Sk&�/�`�D�R�ҟ2Ya螂��
�W�B��	��|�0=��;�0��lh#����Ҩ��J	+�ա�wv��֤-?�~�Q���M�q9�̿���������ꜣz%᳐A򩷾�H��eLY�L*��}�	%�Z-��a�����m�������bp���ߓ
s32�����,x�ۍ쉬�s��&�B���nO�*9���k!,��fDě��O�����.ߩ5`W�f/��n�7o 5+E��)���B��|�h��.��>QPH�����I
t[e�N��y8�&�9{��ݲ�rf"`w�'��k~a����Tr.��P`8�5yɲWg�4f׽�ͨW�!�'��PWgO	������I$����M9~{�S��z�������t��,[M2��bES����pF��� �]�PE�i����A�Se�S1R�؜���\[߳k:]�_�\xH���;KT��V�KY�y�w��t.@�`����Q\wi����Wd�'/�m�wD�	ek� �r�NA(�y`e�<�����!/�ew�g�|��^�m��v!���������L��� �;g�fTX-��K.�2�r�p~=ֿ%��dPKS7��29;�\l:�r۳џ�up��Y>�~Ĳ4�D����+����C��˂�n��FTV��*��@ж��슪�=E�JRQ��=���<,9�?�wД=@8���l+�����G�@6%W*J9[~	��2�)iN&Ri����������_a��*z�FPS�)�_����F��;5i9��p0m�4k��4H�}�{��N�4�^�e]��c;�r U������%�u�ix�,F�2h���W�D�
��І]�V�p�4�.���+ުE3����:��o�LB�:��G� ��A�DJ鈚��#6m��������������hBt�8R��]�=�$�w�_��_Y~�[�vQ���Pe�O/P(�{�y{��5PR�������U��Q�m�{���@QSݮ���x*��-)"�HΞ�����ȗ<�r[$Gm����UuC�z�U�$zr���n4��t�ݎ����������1/���S��#ۧc/�̡_@-��:�v�"��`�Z�NӐ<�vv�iz�Rӻ�ѿu��i>�5���Dꊷ�k���(!���_��x�!�{J-�(���'���ꝲ�@%���Q'�x�\�Z[�1��mڷ(v�/v�].���g�����HƼ�b/��������������d�v.��;��!6�k|Χ։&t���l�d�� �3��,҉����J�_����<3ʩ�c%/jk���c!���Gs���}�^w�s��|���MBVX��M���5�,���YM ٻ�t�����D/ΣDqϫ�{I����B���M͵���ⳟAJ�I�:��S�5����T���}Tt��&./��:�6�yV���������D^C&ϕ����=�����ܡҊ߂��yF8:�U��dc�G��H#_[�x���X�M��f��X
�^J\�a�I��!�h⌡�t�m�R�1���n/�j���YN�5���tQ:���Q�:�J^qr��g�;+������K�_�q�K�SI0	bc� ��r�;��xH�&�K�n�|��}q�T���W�d�����i5�9_�^e�����V��)�`�;J�����%L��J_�j���]���&W��!��Ǌ�����:
�����cKZ6�oZ�kB��uu{�,}���ڤ	�3P[��&H�jZ4��Q�h�NJc��l�!r�������y���9�T�=��{B6�z^�I~�0H�yZQ�����e���@�MSVs�{��n�[�D�>?�9�}���>M��h��w :X����8�@e|��j*]���� �������M�.��~+TU�,���F�8}:.��s��`�����d�Z�A�9��9����"Ę����ߛ�0�@�'5׻�ိF| �W�|����c��[^��D��F�`������9��
�ON�H�ea��$�l�?)�r�3��JFRs��P�>�z\ANt�0w�����us,�ۉ�eO���Q�+�c�y��k��lfF_}��(� -oP��m�H�s� �l�N�aV⥱���%�,����tu�����0C
���9@�?�M�(s�w���\��L�	Б�Krt�?��@��JԳ!Z^U���C�T�@�bI�s0o삠�GbEX��}�BE��2o��m��f��z�� 3���Q<}h�W��@��lZ����Ŭq�G��a=O��:OQ�jS�4p7�	����'ؗ:A�����?<�\�j�j��v�7�w�go�l�"�Y��q3��H���f������c�n3 ��c�KI�a����&$���I#R��{�nݩ�-�f6O�VS�9V��ا�
iJ5��
ʸÍ wH�gY��HUf`W�� #�k�t�!e+
�|����Jʅ�����,�ﱤ�;��s�O�'��}�R���꣏r��miK�w���@	^�~����A�O�Sj��<�*_�r����������{�X�燨��b�L	a7z���G���8Y��"�z��̒�t���]�u��y�O9�}���!D�Q�۽���"�ㆧH#�u2I�\b�(��p ���`8&:h�؊���+�:A�c��2nW#qj�7���"��=T����n�pY��E;������g��ȝZZ勆�_��C��Dຑh���x��O��b�*A� Sw�@�s��ke�IW�Q��r&�S��ߕ�D?�][� Ʌ
��\�# ����T��3��%Y�������i��Eu���F(�?#
�V̳j�\�+���ؤ��d��&���#'G0��U�h��s\��la��E�p��'��7�;p�Q �|C�.���xg=��@��r�ŷՊ2@�+��I;��2�S�<y���0&�)>S�%D����=IE#��#��=3���|[�i�?�]ߕ�<Z�Nu�w�5��ݦHVA!�cp��|��ձ��?�JP��V���x��g�e����49�:���-�`�ԉY�w�Q��ۊ+������S�0>��,��ԧ;@�:٘��v�+����	���řc�&]��nY��z��C��A�gU�r0]�0.�<[��Bk����C�x�����Š8��p�=ɳٝ^��|T`Ӵn��8�v���F�a��չ�7j�F��s��[k�J�|�d��y�GO�fumz��;�3,-2�2P�g	
�Nq�$� �*�걺��_��4%�h������t:�_|����dPC����q�%X��.�p���e��f����g�T�u�u8$��T �5�͈(%�i��o)�8p����[���U�w��ƄL����c��?,]�}p=����h�s�
�=}>*Ir�G	M�똛��^��G��!(P���H������<~)�}�q���V$o�k\��sҿ�Me��<F�g��xmy4�>uxXx���=����^��_"���K�A 4y׳�o!S]8���(�{���x,��Ѻ���jR}00�uҗ��z}{�����T%�raMf+*��<v8-�4x�	!gZdt����B�
�p�CE�/�}�`g��+ ��B҅ZU[�������k{^����h4�5@�G<�]X����0�0.1�7�3��N*��I3
�:>,�Ş�>H1X|��|�['������ۿ���V����⚄�(^c�S]m3�� (�v�^�����Γ�Q�9��677�{rٺ�Ԫa��I�+����l#!>z/��x�L�ԓI�+"�#jQj�T�?�N�n�Ǽ�(�915������ �#��.06o�3���M<;������zX�Q�\��Kе�.��q(�`=�ج�pT���re=�����_U�[L]z1}�M�=QD�{��A���� c ښ̄O ڜ���we���������������59a��򊦺N@t���>P����?~���+[cRn���D��ӥӴ1)e�����G\7;?��f'd[co�>� )�
\絫�2%�kYOG�󠋆�.i{~1�+��: SfC�&v�ʍ�����b�Gu��Ӫ�����⯗��7����粃4��!���MR���|��=�Ko����z�RV���
�3�Gu�C��Pi�u��޴�)��-��]j��i���&���F�������eMw��[Ӻ�<��&�b�4h��*KY��=:���ک�r���&��_�d=|#�>���{��p��I)K�����d�^�ĝ�;���Ў���ݔ���皁�m���-��/��;����������a��c%v������(�ٌ.l�c����Q@%$Zr��U:�!�xLY�kX+�W��^E�h(���vn꿉 F�:|&�J�h�;��ŪO�BS��ygZ��q}����w�5�rt�.ErE�s���-�V�C�۫��6{�W��,�4�~�%^�}�u��b�Ι�m����	gR�_&$i'nʼ
7Y�x�9U����
z���Nb��X��L�޿몑ػ;B�eηa�j��zεD��=��"���yOa.�A�B������S�N4(_r\�N4mH?���t�LI�-���	H��� ��]I��F����Z2W8i>z�������AG��D�;X����g��A&]d'�$���xR6��t����)޸�ɠ�G��㡰�<B�%��q��x��KY搒�`�룭�x��@��-
��!.Ŷ��LQ����eCIV�U�O���V����ð�t� t�ږ�ĺ��+�ʣ��#���q�O���Ğm2������ɋז?k��T��E2�\��3�X�[����7�l1��q�kX�e�>%�G�w�wE�Yvyd�����[����sVb���슕�L��5��
����_+�nG]���S&O}AJ�y9�]��^��L�����!2w{�����Bmλ�{�?hj�����؟�r�v
�������$�\աas��H����~c��uri�ZB�,�G];j~���r�k���������]��L��f�؆�_��'�Rn؂N�ꔱ&�߮Z��.W�\����>
�.��zK/��O,Ǚas1Q��W%s�dCՅ�~&b�x���-�r�)��i<P����t}4���eP�c�ql�Ư~TA{���3�_(��a��p��<(�g񬌤�հ�F��=g�C��Ռm(�[Oh:���O1b�h�Ȉ�B>6m��9�8{���}{�+�t���+�i�f�2&��.���&o�_���x��Z���~��rGvc�$*������B�a���*�T��BCJ���� a# �;�"^V+.�^�T���J^�J^�h��� ��sm<��ڐ�gP�
kD3WA�N^gD���ƨ��������:ሚ���WU�iNb����5����D"��'%��I-�|����!t�Ym@2fPWVF	+��GsW��N���~�}�Q����|}�t��E(��O�2��my���rO�o�b>X/�e֪ &x��R��X�s�ϙ*%�x#v�"�bN���0P������|�O������������]�����bȹՌ&�n4h%����V��6��
m��ϧk\fɑ�v� z���U8�\���R��2��O�f�fa����/^ ��ڊ�Àӵ�Z�����AŌ�uCU��|!�����a���)�
{Br�r�t����t��l���K��dA=������ M�3�?f���լ	�[�����.��)��!��X� �!: �����y�=�s\?sw����x~�)fb��85."����7LdIш(����]����+D���(�x�s:�U{���w}�Xs��~iz"25/_3���]M�����~E�J�{�1��&�4K\ �Š�b��32Ǘݛg[���J�¢���c�ё��f�IR�䵚����S�u�FR`�]�<˱ۘ��� �N>[��vߒ�	/�Ar���>��N�]������;f,�-�+�F�v����׮��D��]4%���L�;�PR�C�༵���P�
�4�o)�m��n~��g�-n�-���߄^�=��$<G�I%�����R�j1�I�!6J�JM>zg7�/]�#J!��ɓ༛S9ѡ����1��3ҜĪc����O�U�jbo�Y�)�M@��n��9�s�m�������2�\�'H����̱�i�ɪ��3�ޠRљ��y{=����-|v��k�[�_����"]ӻ�[�\��t܂T�Fk:K��l,���(fv���G�|��I��m�*�2[�pyQ�����p�X�U�w�nT{KkA�+���kC)놵����5�3(q���0�S�E��u���8uۈl;�2�&GI�?����Q�3�<^��������a�咰�K//�-�^D���r�+҃2���0��RadЀ����R��>!Μ�hf�``�-�U��֔��ע��T>��揕/S� ���ݽ���� ^#^�ɕ%���Ⱦ�c0r�{n�̀Ȭ1���i�Ѽ0��E�M����] ���SGw�59����c9:>��8z��.��.�'K��maz����59�Q��e�u�~��ޜ�J����U(���6���}K���_r�� �t܎��eF�|X���d�f�1չ�8��bי�)]��b6S����~������������cc�_X6kL*�������7�lY;\^OQ�ώ?��?�m�ޣ'�lS"�nT��_�3�4�A��u����?ru(t�-԰� ���\�rgTj��"�S/ fII�q����D!��U�II6D���hK�~-}��~%�z��7Ո2�1 �g?��$4)�i�๒L{7pw	��d���l� ����]�#3~2�W,k~*�~O��k'{��o�mS
�,�M�r��`G(��9�`D�.h]�e���Y.Bw��^ \��U�L��8���EZ��d67�%%}V6� φ&��z[�E�e�����#�d�*U�޺ǃ�k�z�?x]�[2�Y�h��?�LjHu58�d�G5�Qˑeu�:�Bٝy�q��Zh1��M0�+�=��ĸ_���߅�F��̱�}3T1l���OQᎱ�gI1 ����N��6�[w�Z&h#���1���Ʊx�|w��3������6�w](lu�S����k�⫒�{�X���@�8�����a��([!Od��V��MY�� �^}�����1�Ԏa#�u�OS���[�M�'�/A7�勼� N(bZ��+^$�	����g�{K�y��ʳ48��S��*ƙG�co�y����_C<L�`B䥗Gm��J�_߱C��w�/�1~��(]��\��V9Xe���;�t�I`x(��$�Cƅ���ȿ@nc|��=��S�B�tW:8�#k�~�
���xJZ�N%�%�⎔ѭ�T&���=r�
m�i����2<�|��R�=�׋���`(5(k��`fð�<����~��E�I-Ժ  �豊�X��oC�/:b�]�o�1����^.�\==XN�7SB�\�;�dR0vpd_�[A�4i�nJI�%�����h�W�߶�[ �zħ���;Ƹ��ڹF�k��F�rZP�5��.������'@ht�N��o2^�����}���n�:d�����0;���~��y���g�2B5�R��n�Ǧ�Z[�	mȻe��-���q3��(y7�Hv��a�f���Uϩ �g8�lm�A*W�x��m�R��د�Z��}HH�pu�������ʺ��Q&���uD*MvS!�����	ha���>�?
�'�p�԰����� ��UQ_~�j�/�Ի�g�ڳn
�O�j�{rs��(հ��k��'�c��j����y�>��;c����VM]Y���y,01��c�5�wk5�H�/��B��8jq+���b��`�H�$ՠzoi�����#ZtCq!�f������ۓ��
N3Z�zs��u��N+{Xz���r�갴g����~�Km��`휌qO�TxLw'���S-��Q��h���J����(`�>�.���@��?�Z�zb��ɢ|�����-Y?��ZOO�4��3c�Ϭ)@��I,�8b��{�K���9!?>�����&�/�ζ@��^+2�ǰ�R��3���?.�V��9�W��{�8���`�:������Қ�T�8�n�q*�s���cۡڞD���K��� 
�-�%J��T�JYjrD���J�{0�JΫ?��禚;��4a�!��$5Լξ���'�w�~'����rγ9+��'�ݕ�a���WK��^E�c���N���r*�� ���w�%f�$��f)��eUFz	X�Db��<�/8�b|���Sq49���_r�5��W�[�(�)�umQN�O�qU+(�ч*eS�d�x8X�}�:��nƼ��/"����JiW�z6ξ��Wq+C�\aI\(��ɚ�mA��~�l�FQ����ʮ����<˩Z<Y�Q)θ�s�!paR��jr��h�::��wG�һ�w$���4p!3��=�oG� R���a��;�U{���F�d
�u��aE5�.n��o��r�J����aN�ꡫK���!�}�I�,�=�i����w)�k�:mt׽v�E��2�"�C4����dVa����оO���
��qЖ����y{�9��+1���'��谏���d��I�D�Ye�4���q�4D`v:��~l���a�r;i����X�1\��'h����d���	�-���nS��1{�=	6�8vxu�\�?�@�: �G����/_~��k8�h�ET�,����s�B����4�S��_�I���0��WIp���?����%g&M��Ǖ�9��C�RQ<�
�����w@���n�)*�.���k5I�`I�~z��u�۹3J�uW��$�����l�G�;��AUֿ@��R���И�e/��qvq�{u��mWf��B�kg��^%�H>G�Qv�����}����0A�c�%�2PYkA\�����4<Y�<����*��y�"'��-��?�"��װa��u(��A���(<�ͤ�%�^
S�<M곍zO�7SҾ�p�;eڎ���X^�����V.�G���$7p��s�W>��X�-��y��U*ќ��;���٘�^ ���Ӣv���kk�q��d�`��-��z�p����?��ϲͤ�倱�R[w����Z0W�tG8e�����xd@�E�	�0~dB�wM���U�5j	�K��p	&^,P9!T�|�K_��u�穇����}��,����Z��^jc���p��@��v�&��EHn�ўW���rW0=	�8�=]��[��?[k����ҹ��h��?�g2�a�
_M�c<�-eR�|?̅3+��=-�9��U���r�B���M��#3#���w ��,�{�3�f�i{�)���q��Γ�@;���B��'��j��F[ �,7�3�O_��rsJ�#�s����q�ʸ����af�w}JJѺ����|�˗�2#.���C��4��һ�GJ:�iVmi��w9��-�E=�l��I�ځ��13Tp�D�:������#^J,��a~�B4
�&�i�2[�ῇa��K��!kW�Z� PQ60�T}ʨ&�t�����_�&�Hk7�)6���.֝S����O�-��u� Ӵy��*�h9���`ثΩkD kB+]�Ѽ'T�0��@ʹ���#)ГDB(��3�{�
�2l�:*���w�Ss���N�S(X"�)n'�V�[O����^�L�@�����k���H�.�V����9��4?K~ l�gc��a��24�]���-Ή6Z�p��],1�]��W�1�F����\<�������ߦ��ηQ�iˆf\�5>�1`���U�z�M(i���5a$);[I��qC1���n��4+��feoL��c�f��gB���t��h�=�ؾ;Y��+�-A�:��p[�V�.�t�m��X�]i��T-4��>�>�!�5=��A�fE0���L(u<�2��Y���W+
�3a<5[�.��tn��yeIm`����8�Hi�o�).:�ȋX���R�9T&��"Ry,�C�KqF�c�Tg$j��1�	ǎ�@�hK�����_]Zi���ᝠ��!�R����O�G�ӱV*����>���pC�3ȿ�>����cψx��h�]7��3��]�@��C�<�i�G�W�s%ך�xD=\�]��شrFF�p\���2=����-����
Z�E��[�W�.�[➝�&��`{����5��������p��Y%��FT(6���Ȅ�R�U+�X٫�+Ă���u��/ʙ�~���t�
��ᱲ�X2z2<  ��S��p�smq�j�L	�%U�y�6���[��|��`�c����zh��lF&|gp�^��?�"����?s�U�ڹFd\'�Pz��S��B]�{7��l�\�q�m��o"is)c�����A27/�Ʒ�W��MW̌�����/|���u_-ȢØ�)�0�EG)���/db��EF"Ƌ���~`����c�S �({a~��af�Mxo�ɥ�5��Bt��>zg�'_$�[w�Q�K9��|���g)���ʿ)��ᔦ�#��&�4��+���_��ԌyL��^Y�?�gؚV�����3���M� ���D��\KZߟ�=i�D�."z�����ʇ�E�CY�EK_�kyn�u�e���nL���8����)��@�vR��Rf`�O���0Ի�<�
Xϙ{��?�(`:���a��O�!�ymn&�Oh�f�]�Ԓ��J��fKS�
��:�M�u@�"�1�h{i~��29�]�^�6Ƀ��	�
�Nyy��<c+��8Qw�0c��yA�F����ܽD� ���^?�G̷�;�eIYJ���#�T��dkN��cV����-P3��^�kd��m�'b	��Q��%Nv�`�#��`�j������>���$��[ ��o�w#�-i�����G��R���[n�5�Mщ��M_���)?� �G��Ў��'�3��7R�;e'��&5xŎ�(��dn{����3g�j!+�Ui�E	��t#K1��ۡ斮܋�]$Kv�V�z���N
}}�Z��X�7E<L��J�5�)5&)����̷���}�ͭ[j�I�~� �~�����8$�:OB%!�ձ��G߭���6l�{��Q�}���E9��X�s����
�r���@�-��彯�SO�v�j�Q$�m�@�@FE����X�5�_���!���spm�2|>��N���`�ʫ���B�⫒���i~����ln���il�#k�\J~��&��w��mF��5���j�������+1q�/��?;��CIe�VIo%mt��f�o�l�5|˳
^��6qx6���#�Ӷr�>�4�a�G�;=��%cxX���R�w�%�I!r�+��\)�c�h{|�O�����6e�Y`ޚ=��6b�Ꮵ�^<�io�.n�6�H�v�i�}
�R!}�I��6n�h�ǝ��*[g� ��'�BC��LHH��\��?͑/V�Bz��cɋ��<��RO��kzm%�V���պI'V)��^1��J�Z�cEZ���-݃�m����R� �>2�Rh?P�SyU,=��ɸ�V���7\�H�^g��e�篒H�dFE����(3���{ͷ�!]��3)6���V��"���-�|e�q0�L��z#�E�jR<�<�7������9R�©~j
~l�j,���ӻ���W��|�X{ie���72�eQ;ym�"�)� p�d
iWjx�����w�>௅+��I���_3�Vr�`׾�����X��5na>u=\��'�|y��~k�	������Ub����m%텴`��&��:#P*��t��Xլ�x�\��y�>�XH��R�X� ̪�7�X`��%'%S��Umd���&;}=��-Ӽ�KTm��~�'��I��_?�U��C�Df{�K_�A�E��{�c�����$MC+��77q�H�: �_�rk!z,<'���Pޚ��0f*�Ue"�*[��Pr�F�|.��֑.9�F��Q���(c�At����}x	R���B��?��Ip�����,��a��9�ΰ�v!'��O��Z8�����F9�l�ȵ�'��	�OvF�
y��ᨈ��4�<$!�<�~�FNw_�@)�Ȼ�-c}�>����6����`�Mشŀ~�>ukivܹa��Y�"�5z�����TV �+H��L��FC����v�s�?��j>�A������D�L}+�NӤ�9�A��.~U��!���'���S���΃9P-��IQw��ܱO��޾���^e`ak�U��-7`�6j����oT�CJRN���B�g_Q�z���.^!����ʱ��Ք	@/�rU���Đ^�j��|ޥ`ί����@��V�gB��S���ݖg��y�<\3i�)�F߰ū���b
��UL���j�F2����#�z���?f�=�QMNG�u'*#���l!�Y�`/�'�(���W�������IǢ�/?�`>P�k�	l�Z2R+¦&�?f7: �g��a�z�*�@���_.i�%���eŌ%��x���h�<�wa�m_�����):�{(��
#$��H��ax�0f+�H�)�c\�^2ay����mQ>��i�UR��$��-�lĞn��`����eL�N� c�v����o~�lL����n�����d�W�X���|k�v�����S���=)OK��������qСk\�fw��m�>�ɒjS��j��������_�b51Q��y����C�U�а*W������wـjKKE��X'���hf�l:���V_��`�7��4�%�w�����	��y�(�	ar,���0wd�S���z/���>}s��xv�Z��k�`�c|w���4�����/�nb�s�c���^ �$q2�kI���N���$�j]�Rں.��3�E��.�*���&A�'�f�&A~r<��;�
䁺1!�>+# �ǿ�x���Z�$��i��6���kl��BB��OF�� ���X���@���ůF�s(�$��d+jw�_(+�'�������1�+��*��ki!,Ba���Q���_�7���S(�'���O�Rl˹/����㊿����y�y��.H�L�ۿ|Ru/Ů4�m��`pes_#CF��R(yW��t����1�B��z���g�}���P^���	��.qs��Gk����q�Y7���i*�`gV�i�d}M�i�K(��+�!$I}�P�W�rdo7��Ըdn�aS�W�`Oo�[�6��*LA�N~�C0�c�w������GojW���i���� ٩��~�����J��YJ�|�H��RwuZ]뽨v>jGɮ�.�ga�Z�F�wc�d}����Ƙw�fXb�.�T��Ν�z��������T��ͳ��β�nM{B/�$Gg�WZ�7��+5U+b�[&�3=�0��JМ�yo����:#�ڸKw:F�zLLs�_>|����qZ8Db���7�I[ΙQ^���H�&J��%S��,3 Ҏ_�y�N��aJ�-w�4on�|r�=>P�)�*=ָ�nk�h6z7�ɂ4�{V��r|]��2m`;�����eC��U�3�mCK.�����+��Y�z���wױka�S�'�豲IZ�\����rH��d��[��:{�W��.#��f}�����E��|�\l`�:�+�+g�� P�u#DM��ϙ[���3�{�[�\_$D
�5#B��Mb)����ޓh�Y�Q�u��qcA�:�/kJVdF�X��3f�X�G�sT���٪*3�Q����c��XL���N��I� UY�;j�nL7�v�� ���j�*�]\�	e�EK�p:���ǁ˕]	@g��+�ڤ����\���s��&�\N��t�Ӓ�!���}�/(^�g}�$�kP�[4W���>�*nZNX�4�iO�m?��(�Z��|��o�����Ǧ��z4��E�ȥ�n4yC�j�bY��Y}m=kΧ*��9��H��f�^֯�C��_s��YqL�$��.������JMl�e��A��}1�-,���Z�;�k�"_��lʉ5ڗ,G�x�G�?�=�e��ev��d�[�=�	W�Z�����Ս-��k�~��{S��d�]��������Y+�8�;��f�sz��˄����H�]�x�X3i�˼��!o�2�(R��y�98À��]���Z�g����՞�=���5�u�q�W�!�%�S�E��,C���g��n������|aa�NrV2�8?ŏ���l�ĬB��k������������|_{����^�Tv�qpe�ݺ���X٭�(������cכ'��%��#I+�,� O�����x���;��C� i�â��̖mM���_���&�3���_%�ռ�Ӷֻ�E��Q(���"���uc5;�˹gk�m�Y6;Zbc��E�)=�_+����zq�*���B��I7�B���}ޭ.�z�+�5����,�RQ�~v}��C�頌��T���D��=8�v���}�'�'�������u'�;	��g��g%S���1��FK�@	���w�Z�k긹����{���tk�{�Ek����}!���}>�:&�6+g���cɐ�Q�bs��ЧKl����iZ��i�m��G�by�Kie�j(�ۛ�����F	R�!�}rW��@V�������܀�&��4�;`S��z�o�ț�%h�R�%�C3�*R��x.8���VRU�bh��?>��CXa��z(�Vl���R��8ƥ�RBr��}���4^�g�׾ӂ+33%8��8R��W�Š�YO��<l���i���� �y{���7mj+��qa�&:�<���3��Z��Cl��M��\`U__�Gw����&
�O����?ʏ1iQ�-W����vҧ|yݱ�Bp(�v���=/��������K�
��6?C����"�+�-?�x������(A������0�G����L�T�`�{9�[E�k��E{�ؘz��b����Y�g&Z�jst� �L��sٟ�dJvb&��j�h���U�7������KiY��c��:?|��T��5���gf:J��O�g��0ܸ�M!I�6�f���e�{m���q$���(�>��]���&�Hc���V�n�)?�MK���e�Xó��C8��Y#ϻz�M�Zi9>��@u��馜���;@���gk��p��U77�D�5���Y��X�����K�G\3��=]"�W��W]�>3��c��'�^ew�uro�.YA�|�)�&�z"X�E}ֱ:.�SI�Yl��ʆ���iR�a	�\ؘ�P2�%����P#�Nqࡔ������	xc9\F������7^}��
�Y��2[;��ê��""��{.%�K���b�K��D����S��S퐣>>j{�?Tk	�r����!��^���S���������m�|����G����ީ��T��J!���Q�T�殐��~�\��=)���~s���-���l#�\��nX��_�������y>��y��+�I��5�i��H7)����f�a=�9H�5�9�7�;ۖ���[���%Cp�%��$�{?������RS��gˀwǉ���ŧ��`O=ْ����W�e!a�1��_>���Q�s�=�H�m����,
�#2)�L>m�޷��i�P���)L�v͢EG>Yv�(S��ތ~���ͯRl�P�?aדtKp����& ��GR�:c�$�DR����F���ASE�����f ��x����1�)��G7��������pU?�D��ڎ�F ��Q���	��Lے���Q�f����{ҝ=�s^����_x$��2I8��˓���S7��S��UCS6ue�B$�����m��\��>�<�V��ZC͌ݙ��Љ��Y��p�u8�@I���C �P�X�IyD�H��LX��|M�G�W��e%A�_��9��۰�bVd�F�pp�h};+s���]ѥ���~���%�P�1�Y�Q3rݏ��Fа�r��Ɣ�{�k�����,�����=���K�5�����i�M8�3�y ]Πp}�ˢ�ʖ)8|wY���(w�;� oBœ�,��p�E�Y��s��cG� ��y����a|��5�!���G%S��vS��/��K�3(G5c.8	��wQQ�����GMԯJ�<MZ+�����|*�����鴟����'o��G��~���n�8,��o�F���3�RWv�U�=$���`d����#`D]3d�9}�������^jlw�2����ݳ��@�f�̅��� ��V��՛�-f�����m���vc���H��SsC>��ܜ�6�����e�V�,r��H]C�^�v���\y��S
�	��W��\�)=1�_����b����~ί��C��b.����Id���j#":\ 8��(�Dֳ��Gg]-���@C�+O	��9�+���T��0�jT�\/�]Zl�3�["Sh��Ci�>����G֖��w� ��Y"YНJ�������M�Wd��z?�(ڿW�F�?�u���� 6=��2��>���o*�U��V ���Up&f���z�#2�;g�R>�\�/B�!%��{������xv���'�>.,˘�IAq&�'��&8���>��ҙ㡢M�Om�߲�@\ ~}������1�$St���5� {^����r4t����~7BA�����k]�KY���w5�Cg�{`e��/���b�jc4�_��g�xx�o!���~+k���������,�K�?Qʞ�����z+��]���<�Dv>�d�.����v<������g�^Kߚ��J͠r�}����Jj��or��;�{�e~d���t��c�6/
����0�#��Z�]/}1� �n���b�y�z|F��~
�y~P�����*?���!d�� W����˘��U�d8�9�/��P ]P?ς?���X�gG��g]!#/oh=xir��*�%-ze֪�=�gKXv{��|��X��ƹ�;%���#�'�"7���Q}�a�0���������I��\En�C�b!�-Hx�{�_�45tôob�{V)����~T�l��j@Ό,x��k�|�&|�PI:��"W�+�s�4��x��s�R�Dw�F9� Y7���<����>5y�4'�_F#����h���.�
�K�j��U�&�M�vEpx�0�Ey��3��o���C�ö@u���F߄:_Kk���M���Ӿt4|�Y���x�%�|!���<U�P6+(bO��0H�s;m�������ϰ^Z�\Jî��[�3�p~v8$���S�D�na��%\�շ��|�祉S�������9��H�$y��u�/а�����+J�&�M��������Z5����|�ۏq��S���l$ǯ_�������Xz���W�25���۾�~�z�ȗ�U�	P�If�5�*8N�j�,<��PZ�;�ѐaT�Z�C�ٗ慱�O��5�15�kv��L��͂o�<.k@��c§�u��[��7V�tn�p-������̀��6��=ʆK�\���&ŵ@�|�?�;���p(����t(����Y���L��G�<P�v�֚_<��~���@�IX��g: �V���@MJ^���Fi��]���i�
�j$�tn�wCip�.*����/o���w��s6�.��G��`Y,;�.�[����>���p��HҴ�� J����A�9%�9�[U=����|��a���@>�����C�:����~c�z�Cg��E��-S�3�礏��d�g��W8ĆC$�UV��bL�s0V#@	��:�r��;#���1V��;c��曕�����ŽRF	�u�������1�5�SGx�*n*�4���
�&�mc�8��^d}H�3��nb�PB]"(�v��_�w��7�j�_WA?𶨁K�%��#Jѓ�7��/��iϑ4gӡr��/��}e��i�|��%[�H��u>�ߴ,H�HI7iJ�Ti1��]:p�M��0u����~Iޫ��W	�uY�r��p�U�<}*�6�54�Ȕ�����,���9�l��X��,yRNּ��� ������Shl9qqy��y�A� �gw����U��~P͛��*���5j0L�c�N���m��u�\��Q���¤��X�͆��,�vV�����Ti�ӡ��e���n����麪�R��LG��40W���0ճS�s����f�Osw��f�F���ՠg��p�����U�mA*ROo�H�q��ʂ���5�^mrJ�Y.<�I�����������&��x�2%e;�wj�r�0��|�'v�O������̀a�iπ�$�/`���(J����Y�̞�G�R
g��	�����K�~�;��M�V��)��3U/��`m��O�ID퇰wz���ˋ^���XzQ�X� }�#���$��b�!�L��/�C�F@ȯ�'M"��� ��Qm���g����Ņ��,��� ً ��XT�\��g�9v`40 ��{��No�+����"���Mq�PХ�7Xd2d���'�zT�-jb��"i����3�8D�<�̼�ہ3���8San��]����D}�oۨ�:QQ��e�e���n���?�-5�٪¤o#�*,���/<ߍ�)p��z����O{����x�
�{�4A�M�⇍�erijA�Fw`Z�٭�����)���S��#I�z�1�Y�ZEކv����X��/j����o �s����I�����kP�ە�moܶ�6��r�WI?^[�7x�,նZ�X��yR']�3;%���;"Z~���B]��ُ;S�WC�*�l:�ۘ]�6�}�����]�K��CU�hN0�{W�ׁ�I��c�j��׬����k�bQN�v�ڹ��Gט�O~��Q���?�@��X0�c�.����Y6 h,l��)�m��.,����U`	Z�:��i~s��ǳ�@S�T=�+�(�@��|�!;ٮԁ�����r�*�WT�l����R6sMS��y���1�^�?E옡c}F���/�����?��(��A�/¾:�[a����0��HRER3��l}���@y`H�c4����o\&�Y/[_������0�J~Ϝ���?hq�6�����ݫeW/w��km��"���Qu�k�t!���dc@FBa�is�X��4:0P�:s5��b�#��#.��J����A3�o
��b��τ�3:�'���H��o�����妁����v́����w�&��:��l��� ��/��V��Q���'�A���Q���k�M(�ZV���gu��w+�n�Cz/��#��E<�G��{�f/|��%-�2�lb���s�
��h���Nc��3�dPV��JXئ�d������zvmFj��^�9�H�W>&=�;�'ha�R2[P,����P��n��p�E�8؍(^�?%��w������K�=8(rd��<I�8�buX���x�=g��Z�������1]���M�rH��F���
YGw��b�
�<#r�4.�(�[׷^��5�49J?�F�.4(m���JZ�;��5�6�j�Z��l���J(yQ�^�䷁u|�M��{(�J�����*,�p�kQ��an���� �mXy��{yZ.��K�$�,�yaof<�g8m�T�;M����<�����3s�5W^32j��~i���)�D�u��y�*oi�6#�ހ���b3�}�WYv.�����B�o���-�B�j��Z)��;SuI߈g>����s���gl�Pf��>y�E.C(�TMX�_+�Zq&�qe%�c��//��5����7Ly#fO��G�n4;�u�?���.-zu� �ZQ�/������Uܸ�]�]ohW��9�f!�r�"7����ޥ?z�������Y9���E�t�q�I�s\�N
�i�B)-;����5�6�gR ���׽2KOD��x?6�X�Q9�|DΠ�y���ѭ��>��`|\q�)Ԁu>o.QI�eRB�g��C���I�A��1�@�l4�����__�a/e��}r�O\�a�A�����B�Ko6(T�s�y�7�m�x�Xm<���=�۹���1��h*�Zɧ��Oz�ީ��I�a�c���ΰ�~�����g\��|O����*����ƒ��O�Q���MB�T&�0�&b�x�Z��Đ��o�]���$��$l<e����{7_��a��g�����c��IXQ�VK��_�֫3"<�~RLË��?wx_�o��K\]`�����yH˽'�#}���W4����>{�@�L�}�cJ�Ӷ�a�!\Q��;"	㍺��#ww̛I)���<��M}�:�>�7����*�j�'��hu5�/�L��N�sԅt=zy�>l����SK��3�[�R�N��JL]�u Al̾��9	��<M��-m�`S_��N[T��oT�sى5����sMiߪ� ��n�\�4�����������Y��݃6�|~��?���0���$���<.v~�̒g��k�.��o}+R}�(1�Ml?�k�t�)��H!͝K�7�������Q��ns&��ِ�\�(Fw�T�e���ŀ�Rv(Vɂˉg�J%�7.f�wm]^ڴv3^�a O�|G�p6]�m��}YX��o��#��h�x��,M���Fh-
4�#_�}A#ǰ�5��o�2�_T?�}�>����<�Ħڹ�����ޣ�jQ_^@uЕ����bi��{�s����9e�p��#���,�.�oq1ٍ����9-���)�e����
�,��o m�.�&�(_(P�����(ƶYxӑ3�+Hœ��/�
1�!d3f������Žȣ<��m�xz����k�zʬ��~�V<�d>�H� ����8h`V���}��b�V�n۩����]R|�hB��f��(�菧CX��������=]��JO���pi[���6�ڑ�Ae�,�攮�H��?ϝ՛�9p�\�Y��딉��~���NMa��\�R�+z3�]H�8��o���f�*��k����}�*�Kީ��g?��[��l�-E�(3�u6.l���$$��L�~����2�g{C�7k+�=G^�9�۠t��F��<�n4�K�̈�0��n:���YOn	��)ˋvɅ88A�g,X(1oF�o�c����}��#I'?�ѾYr�}v$��4l'���M��\�⭘ ��	���
�ς�n�P}E��Ú�ȱrkʦ�t��klر���9�a)p��h�[q�'Ԡ5���( pK�Fq鋶 ���o@���e8��fZ�\�D�_jU)k���+h�@���4�G��+j����H�K� d��}�]�!L�׊s�ư�ƨ �rbX�D؀"x�|C���������Sz;�XU�c���<��`�����q0�.E9}CD���[4�z�ػ񄹾�c�����7qm�͒�	"'6e�B?��8�4�T,��D\6B�e��P�I��h��E����\�JJ*hRӴ��^��~�ǚ�����n55{nÎu�������G�;@�i@A[rs[�;�����#�FP��2)��ܿ�z�!�d��=���Ή3X��lo�UKzs�(}1��̈́�?��F��
�H�'E���l6�x���\K��.���*�Y,^�u���6)���y��8�R�`v��MΑ���A0XǕU��\���x^)�,�B�ajOn4&�vռ��0-A�5��2��)t�ꨬ~'!��)��5N��඗�N�Civ��qG�w#_{�QF���"K_�^��%�[�\�Ŷ���:3�)ʕnw�b׃�f��^���Ы��Yy�گ�E=KuIp��Z�w�Y�#���|�1�����/?reF�>�r�a&ՉԢBH�-)Դ��)��G�	�7���j��{��Е�p1��t@L��4�GjlaW����-��i��GI#��wx+�.�UWCt��c���ocS�z��Sם`�
�H�z2|��:�7��} �XS�d!���,e]|�۴V����+������������m���kgl�i37���Jo�;鲵��h����Ӕ>@�@憐%߱�j���Z������@�jH���9�Z`y$)D��)�&�sMRt�񒽮���7lX�<���N:���2:!ݭ���_��;�r�v��|1��C!�O�
3�i�u'Ĭ��۱�t�*O�Vy��Kg,��i��d��q-��Sm	��^V�T�S�o-��z��"�5)J�܁�!�ʹ��Vq�(|�]c�Û����b�68Z6Ĩ�Ǽ�CvԘEk�Օ��F���*��~�⠤�
3���ţ�����
r�'OU��PQu&�ݘ	V~�U��]��n���Vy�d�:�3�6%�*`�i! Ƒ�������%E�DuU>*�*&,U:��)	)r�Vw(�����o������ם4�2a�T�&{�:Cz�_#�sF7�)[����k��.�N�����0[����.��4�{�m����5�<6�X��:�(�
���ІV����f����JO�`Vv��H
��K+t��r0�xo,+�gC��[TyT7<�υ!�s���.�o�TId,Pbr�x�l�\a��Z"5T|���� ��q�ꅳ,��zN~��f�ך�-T$U:x�;8}�"`&%bɟQ����X�-�M��\~�t��j|0-B�IՀ5(t��'�N�C��ˡ���>}a6���dc�|O�0<0�z��W�W&aS��0���H��A���� �. %!��)�ҟ�#�v��#��U����Z�LL������8�OG���M��32tY�\YS�N��H���'���hk:�
ąN�i�Ƹm�"6N^D��?�Je�G�Z� F�T�`�| _G��$��gV��l4^�̎��+�3Q���q�mG�iV�3�',�N��v7�U�N��Y߇�ʂW���O��G��U騁G�*���~ܳ�G��G�����ɔ�HmC(eK�smU֥��?��	\Q�4�1c!�kʭ
?o�_Y�9�J�LF�s��.��v\���t��.�>�X����o]G�l��i���f�l���Y��&��ֹ��\ς�إ#O���?;�+�/��^�=��T��ض��|XA���ݔ�fY1d�q�ɯ''-]my��g>�H|�5Q��`d\�[�����9M��4)#����C�Ǡ��^�%�/fa~�Ob�b������I�\�����G8�Wn[3w�w�<�1	�S�M�hE��p�\n����H6i�,������I�E�-c(�I�pC@EO�Ȣ�����]�<�n�zFQa�h2�������[���'�H��.*.)Q�|�c�����ZZ�38�s$�o�\�ѩ�݄�����!,xt���I�bP�-Wf����	��"_�R�/Mv7W�.FٻcR����g��_߹i}�-�:�ͫx�t��E�)ϟ���-X�mI��	��G�b�EČۤ2���@/����ث�ɂ(�Ц���V"�S�`�[�0�ͣ'��]Խ,߆�(o��"�a��l� ԥL��jޮ��8�e�B�aw�}��ެ�f��,�뽌;�i��U/9k�����场��Q/@�ja�_�����QK�-�o�Fv)�$��F\�z���s�|1�B�F�0�$4���}E�W�i#�U�P�A,=���BS�x5󌺃��C���S]8���� ���Jթ33����h�yī�9X�E⦙�k�3b��t�o5�Q�p�Ї�t���!up���&�2�z�/�tUd���g-�X�����c��B"����sܫb�y
A�z�%��Zݻ�H��Y�v�����F�lj�&#�^��h�l��/{@��-B=+|��tu�S�h��u�\؆���b>Z��̾�f�e���j�^�ѧ�^��-φ;�(˴_�q�����&{y�����c���CWMmM�>b�3c�n9 ��!���meo[,V�ğ�7��i���\^��I� ���>�W+��W�&�_:pd�x2�0�����ӷOY�U�}�T���[+p�d��5V`�	�À"Ç*��1��g�"K���'�N��2Ϩ�������|��i��g�]�� a���g��:�a��)l�L�χ�͞" X��h�ų��J�!��ѝ����q>�_�5�O�>�E�/�X1
-�0���%�7���}����4���Q�9fT
��٪�4�i`�����f�N��Jˑ���'� d��Dyu�P��y�X^�����⨧��G���A��<�'8�����{�/��R[�N-�ڻt��:}�%@��ty��O^�;�,�y�>{�=�;�]+Z�l�E1<�J���
���h�G��dOԈ��`?@YU��I��O^�v a�'���K��_����QW���09;;�o��wn�R]Ò��u�)��h_���y��E������CF�yyk!�g����(�>X�;}at���H´XMk +�ٹ�0lGv�La1�8���d$i%�OW�K
��+/�+�ڝ1�q�/����8���<�Ɉ^{լ��� b��&G�Y~���_�x�������E�$�Z���@4�ه�-�~#�Y#h��!n�J���p�Y6��D1e)�zV�
!N�`j�����rʛ��e�u]�Ml����?����aY|M��'�Á��)T?���r��L�g7 �����kp�{B[ME�Cw��s�6ILҝ[���Zp:�8�<�D�=�}>��'s�ہ��NO�)k���K���7
o���@'
E���*����$S�{G@m���E�Z\�B���}U�v�i���m�cS� �8�3�8�?[�j��L�	8�0����\�ޑ8�O�V��+s�|���v�z�	�rZRٕ�:	��
Bo��h��z�s���9��Q>*�j�^~���ȁ풗����y� �b:,���r;����'"����[Mz������Z�VUTn���"�����)�����E�������p�:�ہۑ������@+.��:a|Z��ɧ	z'���ӣ|��l��.�ށӍ���hTd �����̺Y7��i�!�皫�l���b��?�Q�=~��j���7y�f���q�	�a���wf�FR~�m*0���|z��:})�{wR<���nЖ�(Ds�Ǔ��u��}j�̂�)�7w}IQ��ζx5Q�nu��`�c���(��P.>$�F�x��{�5r��8��k9��,LOR������-�o�I���8��_˩�d|���i�q�V�`���.� Z#���o��=�G�D^�"�^�Y�ϯ�݅�NI����@ٞД��.��L63 i&d8~�� �(�bD1��H���+W敧�Cj�Mf�`ٕR�y����R�s�e�-�_��Fw��f"	#����y�5��� � ���˛̻[&���dd������Gr��c~��	�)6�TT�P�S��&�Г�eKU�QqɃ-΢�n�jg3��Ed�w�x��s��|h�S��ٷ>$�0쑈+�ч��^AyG��(���(��z�+ШJ���q|��JW��`�N�m��D�t���2{��4��jdR�Z2�<w_3�s��ad�=$��BVa�mp�1��k؆`H����N6�f�{����k�ߦ��������b�q|��I��-yA��%,����0,$c�_8�6��A�7�2����d3�X�g��Bݫ�z�F��Y�Db��2u|6��>�ҫŒ~i�J�8�bf���e������~��A���o�r�q��A��-�6G^=�4��M�)9&r\�\+�%ϋ��G=C&�ey�D�11��{�����.³��jo����L�I��l^0*��k'�������!Y�Oh�^�<#�?�2Ԍ�#|��z����׿L��v{�w��N�&~���\L�?@��73袤�V�_��|('#��$������i����^/MdÜͮ�n�+�<�}���"��۩�>�E���6hv��{�?������ci3�D�b����+�^�E�5�k��5�E���s4�a�xx�n�j�c�I{�a(�;�&�7��L�B#�3����
z�ц9��6ռ^B{ $n��\�����ؼ���XD��1kyo�����Y>����l��%�wfL"�P%#Ѕ�2�e�7} ֱ�6�(���2��6t���u{��q�=���`}>�mmh�#�b!1�
.���#t����Q��Eg���o���oլ��zy�k=��<�d-�F=o^ۈ������W�s{��<J���<`!�cmL붦<�G,��=Z����F�ߤL�
,}�"�(����YO]�@5[^�f��xݴW'O�W>*j��[�e��L�;�-�_�?�[�:����7!�C��y��b��� ��`ؗ�H.ZNp��]~���n�^��D��������.�~��!�[�k�!�>��ۑ4����k��`K�v�Vv,0,�R��TAq���D2��0y4ɸ��}���Ge<'f�����h]� �[fD�{��`�\9��e��>P�2�g�n���/�0f�����2��~����j�w��8K�y����|��MyޠTٰ���|t�97�>��AT :e�7�8韕}ѥ� 9A��\~���m�I׫eɼ��"�_ƉP�����	�Ǯ��B��5i��r/����3�C`�TyP=2��.ƄIG���і;MG��=�/X���&�?�7g�6�a��8iô�슔&~���]�����T=�ׯg_����}�e>�r�"����w9���=�-i�g��z��V&M|:���NZm�����3�_:���P�Ïs�����̐�\�<�gi�Q���1��\���Z����o��1�'�A^@d���w�6kX�5+&�?�1���哣�m1.�=b��P����duʖijfa�w�ܽ�b.��s��Z3�����zd��c����*�,>��?ƕ�p�{@�A�~ɋ�)�׿�h%#�f��sԃ�.A�=�
�x?$�g�H����w�Ա0���	1���а>���/���.�+�k��[T5r�⧮�C���5��#oXX��i�����W���6�Y���T��7�^Wch���'�,�_��ZPo�����Kp�T�V���)��;
��7���i��\�5�eTG_�X2g�I[�)N�ƛ,�m��+�>z��B"d�A�D*�L�I�6�vWZf�������3V�P~��Ҫm_/1h_N״��>�6�/Jճ]�Ȱ�0ׯ��W��'�l�g� O��>��;��6�~�'%���S�c�q/�W���zfO�Y߰�����{�bf �Nތ}T<"�LY�H���{�qj@f�j���,�p���PT*�w��o�%U+,����U�H�r��Hod8�'D�G�6B�9��T���(��F��y6�=���UZ��Tl�@������x�e>vuQ��L�Vǔg��I����z�E߼8�U��ݐ:Zhʰ������P�I]����:X:D�@�Ї9nL��@2�蜰�<c���gNy���:��1ň8�ƛp7�q�9}8�w}VnF�F�}~~U�>��9���-� �b<?O�d����}��t�WS� -�5�.�-��uT���CF��`��������d�J"I!xJyYM�}�&���Gyy�;�l�"�e�p_"֋���S�Δ��H�������m,�u��F�U�~�� ��I`l8G��(��d&� �ci�8��9�5sT���X�tJ��$،y��;���S-i��z5X_��H�����,1	G^��@3~7��K���~����@.�f�;��f@
��ÍvF�]��ZyM�j�OR� �u�v�-����4"�noo'��O��rC ��*a�Vo4��^������$so9�����l����|��핁�M��
�d)?��Hn�֞����UwU�����!,i�C@�'��E���#�&�Kv�k��,�_o�5�~��y�Vy&;S#�f��n^X���U�j�C����%ԄQFs���[�+�߬�Ton}�����E����/7�Zy���Z;�[��Ȣ��1F'	��:.Sy�Ő��	��M;�"�u����m=0ҡ��Ƙ�9?����U���6������������3^:��u�8װ���oVb����4�>�qYw4}i(�Ӽ�B��l�r%ɚ��`����rH~��,�#�^�F E껬怟��Ƿ�H��a���|O�����]�k��?M(@6�!�Y��}Ø��Cr�ד�@Xo�zO�'��ߎ��Q�7��p����
y����.{��%.j���q87��1C�f���\�����D�.߃qUt1( �Քc����/qL���l��������-ہ�zY��Vj�ؤ��û�b��!�^8���ƂE�}/!v�"Ht���bg�yQ��f�}]5�})	�iIˉ��7k���
_�N_7�}o/�SG��/u�M�)�b4��tw�3������A�>��xt��J�T+�RR�P���@��+gR^�n�
��X�3S՛~8�z�"B�qUD�������֭�o����m�O�������@7n1v?N�;�Eդ��`�k%�\Ύ��P�u|#�t�Fԕ����T�c�W��2-u�B,���d � ��g�e4��#RK�����+��v�e���>9ha�E��2�w���s�����6[����yu�"r�
ޕ�4������zYF��Rj�|t�'��{��iz)��s��i��k�G��f˞4�ܿ�tz�v�LH�flTX���^麪�g��w��d eҶ��������V�sffߪ2��/�����_���{�V��U!�tF�*\�e>9���d*8��,V��y��T�~Ne:�63��˹\�.��P�?�m�LOU�+ab-H	�ٯ��~�ץ(p��4��4�h2ҾAy,�{�g����߿1��i�9Q�:���^�[�y����;�_�[z���E/!x�2��8)�vq�QT���D�t�iY>��GIZK,�8�1��7?E ��JC-�����r��{��ȍ(eE�|
o��*��&b�ju�-���Ŧ��-8�����! �����>ք�nk�F�'��7��3�-s�.�+(H.��3�Z����攎�������9^uM�!�����9������m�L��SE�u�*�]�&td�(|G%J����W~`�Q�s5T�w�8[<��hX/';�S����QSՈ	�_���8�n�G�O��X��5�V�XC�����LvT�tM�;��^F��#e:�[X{�������Uճ*I¶����Fӈ2ZHUB���7����P�m�ʷ�\����As�t���!0��(���s���s3Ȓ�Ҥ��:��T�#�j��3��m�g��?@����ʙ���B6�!��Y����G�܍�Dq�G�R�K���2g��H�S��ݞv+u|&�RlIĔv��ܷd��fS�:�{R�H�}0qd���-�w}t� ��N�yv�6�ᑆc������[���0��'�'��O��"5�����b�Ur/H٬~���^��������O���kf=���rwkv^,��(mt�Xӑ+�[ݾ*s^�^P����%��W�Aa{Z\����KAl4ǟ�И�y^�-�呕�"��j�N�Z�Ot+G�vw��tVs�����~��P��ڨ@����^y�m�G�_����~~�x]��q��Q�����<��|o\�V}wܗ��f7�q��e�(��ؖ��q����틿��jG֊T�Z�P�XK.�� Tdd�z�^p6�߈��j������m�B�������ϘZ����o�D߫¨��O��L��~�+��p^:��]�哎���Y�l��Ƣ��^�ڻʳ@�ꣂ^�e��+qB(e9`�Av��b����t~��c��	�w��ՙ�0�"����,�b�V˔"����#����w/�$G���Yy�>(��f�.�Q#&պ��+�-�����aԳ�w0��:����U@C�,|�X+N�D���쇆��	Ѣx���*���p����;FL�2(�ʡ������������������wT�̗��}�F�p ����k��h�}�ػ	y�0�TʔK�� zofN���7
"`�ݿ^ׇ���+$��d.���Xk����:�*���4�j���I�;���ּ
����@<������E�w!S}�a�G��L����C�!*�!�w�"�^eً.���Px���h �f�qk�t)�U�K�9���ܔ*�t�t�m�#/jRਕ�c�s��Ё�1ȡ�%px�vis�Bc��q��9{C�wk�ET�����a)�ᶵh�r෣������"��nP�V�\~9�H������S�W߰n�'B��I��.b��O�}x�s�g?PD�����MU���m���*̭v֛o�����ҟ�#�û�¸�&�/����Ʃ�X�� ꪰY�J�b���9pŅ�uu�iZt�p�h�;��n��Z�IҚ��^��W/���i�\�]�����G�
�+�E�'ϸ�
�,�B �>��vV��Y�[��I�_�E	�t:߼Q��kv;����l
�t������~:�By�Wkt�G���Cb[�"C�$}�{��A���9AH*�
���ܚ\A9��TV�TY��n�_��w��p�ݫ`R@�x3Fڙ�~]�?�v���bK���0�ɓ�z5�2�d%yN"Z�ea�DJ�7�:
�O=4R����]=N�+N��5�tS�m5л6~,ͨ�����.!U+�"3^?<N��	s���~��$���7�s,��?(�1��4e�?�}_�K�<:���@�U�k؜d�\�����몂[ˈ��"Oy<�C/�N��M��t�u�k3>LP����M֭yK�bHy�i��L�m�,�D������ʃ3�S3��$$֧��v�&6��r�L�8�u�͛���Nw^%�>49����{V}��)̞�)=�8�~�nA�ЭR��`�{�	���/��XC�}�Lg�q߲�G1'f���K��G^���[Z2���UN�����C)~+���Q��ί��)��'/�$/G�["jL�mk�d���=���/�:��/u;��V�n�D�8�{���H��W�~��8�9'~cE.ր�[cw�EA���{̛� �s��5T�$�����5��L/����]�ø�y'-C(I��=���{�ʢ���Z)�_�Gn����h6�'���xI++�f����9���7e�*¶Z����y`�_�~���܈B���	Y_��r�-���c.��L�|��I�Ϗ<q�`:�(g�g���"oٲ7z@��2��������Us��.޺��,�i����b�˅n��5�Uغ�3f��;!�
���!�L�+�O2��: )vY�h��bW��G�_S�g~�t�,��&�߼�%No|ѫ������$���K�B]��خRw�1����Ni�3���1�g�{�ѢtЪ<���R1�-�h]Ų�����!�ȴN��_��}71�/T��ki[d<�j��1c|�o�[��k������zŝ���V��wҜO��y.�H����Mu<x���e��h��S1��\�wXz�c���૛�F)�fL:�}8�k/k�ڹ ���IM8�Qf��`�����1�Ega�L�@��^��h(�ך"uU�!��y�wH?_\3�����z��#�֤��c�w�ic1�<��K����
Ҷ��wШ%�0���[��Ŷ�������-K+�L�<�a�p�iC}���t@�!h�N?0�r֣�B�R��gS�>��~�a��]W5oΖ�tݡ�^u��}�Þ��%�����$��$!��U&B�'�'B8Mݜ�&:�1���2�9�xUr�(�\:�����ֵ�����.�к�z;�Y�C����2� �A�� =V5�`��Ax�ގ���6���[�R�W���}��$nJ��fҢs��a���C*�22��VJ�\�Ģ���Fq-�v�l���sSJ���;��F���P�����N��fG��xe�����6�tzeNS�1�;T�Ê�S5��Hsň�o}�������Q����L�[&db4{�B7MH��s��nC���d1��LD�m�ɡ�F�a�v�D����&����H9������l��X�\�Gd9{��d���N�Y���
dO}�Dul�>�Q)����>��ț�#��
��G>����\ӻ3`\�`�}��d<�Nݣ�-˕g�1�Џ�%!B#��2���po���S_�����iE�B�")BH�Vٲgߩƾ��$k�J�lEȞu0ƈ2d����33��1��~�?p��9���s]��~.3��D�&�z�"��7��^MW�,�s�Ƞ����Hڢ�~��ynqH�q������9^Q�RP�|���ܤ!��f���{3#�MZN��s4��,��
6+�	!y���'߉� \QŐB��0_
��;�#2^�GON�a!����O~�[�B?.�J},��t ]�`^�5$�l"��� �(���$N��+ZE��vد-��]E�;�~\��f�rz��zq����R�B�?ָ+��r@&�����ٔ���9��W��:i���}@T���1Y��z[�B�,*�Jh����S.
�e����"?7��+۔�!�@�f��������7<�N� �+��è��x�*�q�����-����ņ��Jʽ�Eʧ�R���'����O��B�=V惵��Y��_?�f�����?��Z�����x�-L��#l�IN�T�7�8��'�?��G[�u���i
�tOQ{b�w.?y��v���XU�}����F�j+V�K��v�M���!_�
��*�[�֥���Š@��������C!WFbWζ�z���$]a�w������1������I��ȃ؝�$0�J�;WlXi�@|o�����J48uH rH`D�^Z�zf�����&��:o�r$x�z���.��m��W�C<��{��SS�۝� i��Q�U�v��j���bn�;:J���Wg�F%�`��9��t����D��5��)D���\?f��#m?,"`CNw ����0���8ه^�p��=�;}��}�}�Uy�q1E}���u���@_Z�P�'E�L���� �k���w%o���w��AO/�S0��
���چu
%�`p�:�~~՚�#��ʤ�3~V�W���ћ�
�k��Z �_�� �q~�� ��y�J6���.�፟�o�HY��j���_Y.�k�V~����3.�^��7!���Ni������$%�u���&��_��Wu�����8������=�\��%-�9]����Wq8���R܍��+����ɛ�ogp#���VdU���|���:Bi���j
�>4Z|�lA� nt�f�Ƽ^p�Ǧ˝���!�ߕ>�$�%к
l<=�������6�b1@\��Η�3M����c�6�[t�$�m"y�������E~�����u�������M�+�Q�.�0����͇��8�&@�;������cyM��(X8�����"u'w�AI�b"��B�:a�;�Yb�q��"D� a)�C�q�g���S-|镇}{��ч1�E)Zcz*J��0"g֝�=��}�MG������S��g��9q��X�����O�)����4��4&RKLe����^����%U�G"�[���#���[�tZ:ۅ�5������G_�:wPF0�Җnd�%�Ts�mJy�;ߑ��F�P��tY��bb|r$�*�!�[�'������f��������;���˟��A�h(��U�����&�rg�
�ރ4y?�K3h�-��K�vr�p|�Ӈ=�!�f�����G�ʞ��i���Xpı�ۼأ��<���<�x�-{�1���I��җ��V�G��|4<�k�5���R]m��GԱ W�ښ�c5Rf�SkӒG������'}�ըt{����7s��mj����[ٻ.�s�s�z�լW�D��$�fS4�c���e���7�?"0�^��S:��K��KgT��<(Q�M�{��`�Ah���I"���i }?bmT�a��|�٪�Pn�S���!�����6���@p��i"��݉�
-�&Ah&��\!)�4���N�>"�tcz��L������ݩ ���"�5�6�.���x�w�P,eʑ�舄�
��7���e��~E�֥t�V�s��ܥΆy$�x�<ّ_��6��j���̮��ёh �)�$��Lf�Q�����.@;DC�>̗9��Uƅm�&�H��gV�	�^�b�0��o-�w��1�XO}K�^�h9�,MҩE�����BZm�͇��w���V� E*����97Yҳ���l1�%PC� <�lV��Bz�����޵��5v]2��#<=�&�^Lgo��V.y�=cx(J�Br��G�JD�ԝC19�R��������ƿH_9��[�;����A��,�r�Ɂ�����Q������$~�Xyq�]��������[�U��Y�+���M!�Iުs,�z4zZ�8ǲ��o�
�Ga#5*���eP$��.]�$bu(�+�>���݌\l)�y�a~��]����[նH�w��R)i`TkQ�ZBm�A��`�js�2毬�yf�]ᾖ��}R2$��Oٗ���ad=L�lE>{;gR%�H�%�L!"��C���:!� k��:�>���AۑL���]Y~���i��O�+\����"FrF�97� ,�+K��bь�|�Y:���,��r:�I��¤Kᴢ��횇ֿ��Ǐq�E)R�������6�E�ma�fҜfvV��ћ怒�V�َ�iTG�o���R�<�EoA��kr��ブJ�:�y�(��\�����l��#_ 9w���r슚V��kA��Lt���6�f�aG=E��V�lZom��D����&`ap�!��;����Ʃ�b
�p)�H�v�A��N��&qp�f��ʬ�Uo}Jצ "���k����Ph�H�e�y� *!��NȺ`uU���Ԟ�s��gΕ�b`�a��(:��Kd�_�#�OxH�-���������L@��)4�ɇ��Ugq��e�5��m���%�x�$w�&N�����6��y��}v��T�H&X� KEmY�?�TpeF�4zk}�f�
?D�����غ�ɫ����0P��!3PE�Eiw��5�����4���?߀����q�����H� 𬍵��]�8��
;T�����@�0�rɔ{��z���kN9��jDۣE�/�d__��S���_ߛ����N�ͫ=�D-�k�A�ɇ����'��`�C�ڳ~�?V���e�3����7���fr���!e:�Ӿ�����|�	���"��?�g.� Y���OU����q�/9a�cABD��SĊ�}��_k��~�O��f��k��o��t-�_��-���N�jh�'�����sK��"kCt	�[MV -h��`��![%���zHɨ+M��X@V(t5Yت�吓�=*b��ǜ��1��d�yGm� ]�0�Fx��2��S���M�8����'����8M���ݡ���A�_j��m<����q�g�<��0?;�q�^��M_�Q=/mQ*r�v-�/�B��T��i1��r�l�����bd�uT��S�R��z`������5�׫?Cں�x��ykl
�@|��ڎ��j"��7I��CɶOt�|X���l7qKj!�4D��SI�w^��MV����nh!��� ��_�=�4�粰�bmGrٿ�$�˰�D�ȶ%����td5�8������f0��)����O���շ�n�sR9�b����Q-"�v��t�P��6s�9w!B���H����I�(!D��r�?:yȒ�땥��TV�0��Pg���+�u�\�C�y���ˁP�n���G���	�����L���x����6�2R�<�}��ڗT׺�'e�}
��nײ<��Tx�o���LtGs(d��X�5�NuV`����Q���gP��̺X)[�3��\��yG���!�{����q��şÐn�[W_-ZF�n�B��`/�/�C�ݾ��`��`� �s����7	3�r�~��/���g��LFR���/kB&0�I���s׾7 ���+����{(�7>����8�/�h��ѵ���b��=��p�>@�E�����{S.oI��Qŵw}�m^alR�A����!ow����T�q@�����zZj�+�m��E�I�[��y��(��c~����P
�Ud�h���tq	�����$/L9�~6d�����T|��5v�hQv�jk��٨w��YV�
��,?�z�TM[a���w�b6C-�J_��ubLܪ��g��b6"�\	r?Fͺ6�ua������F� N'�1�f�3��z�f���@�t���*jO�k{��Vs`;��U��Οk?�u���n�"c�D�	�,w��"�H��w�$4>	a�f �Hjd�����; {%b_��)�g�'L�-m^��	qa1�%bN���(�vV����8w��b�~PA��@��y��#ˡ���~(��2��g ��L0�/�ܛ�Kk�Et����>�ˬ�E7#�5ǟ�y48�!�}�\y����MOF��@ٰ*�s)9��5�d����:��H�Gl�=��/ɦ+���w{ �GB�vV�۾>��z�M��b	��z��C^��)T�Z������|2��懺Pu\s�uG�[�]w���4ۑEW:Tz c:�.���)@G�k̞wdU�V5�:�|�Ek���XrO�&��N!P�*��^�jm��K��'Ϗ{����%Q���B���X�\h�������f��1���*���e_C���a��ޮ�����f z�Ǻ��C"���{���-�@�fs��FIZ��/����C����_.������Q6��&|���t�������"H�p����86�BZ��}#���)[��G��`�1��Qa��u�G�#�;��ON�$�!��}ɽ1G��4\���r��V�+�6~8��IC�wӋs_l�Gb>�K���J��7#�Φ�GzHR����r�!��{�4�2�XLcD�C�B��f�v��BC8��Ї@CP`���}�v7��ESt4��G�g.�)L�/���`�u�9,*F��@�j۵��a%�R[��i��!�� ����	`ѶuL����U"�q0�o	2�ǯoT�������n.�vK�AHL�ɦ�*�˴>{0���&�H�K�?�(�}�Ü��)+F����a9*cq�,&��6���GC������$GzY��>�I��A�=T}!���^��i�B�IJ����F��C/��j0sVŤuS�Ei�T�Ŷ�O���ꩈ�(�w;`6y0��_|�Г��.z�l�l��y�<���>�0��k�	m5͗���OE�U��J��X�ۇ$i�y;{cJXV$�Z{X$�����h�:s�P9�Q7q�k�-�'A|��?�'p�򈆫�b�xB/�Ŗ��:�քw�3m��q��"A'8]>{B?��LΪ��0�	k���E�|P&���p\��݄Ȼ�3H�3X5��|�y��_�M�#�ʛ/�O�T£����3����� ����d�]fVIx�{˙SgB�/):���kq�W���V�n�@QP�aLU!��U;��6:CÑ��r����}0�7jIt�жx>��B��'���|`s��������@�C�ڇ�Ԗ���έHC�^��A��7���šI_���K)�{_I�^�mٶX��gT"H�gtG�]H�xv��G&�o,���"�:��s(��v���ե<V*ou�%����2��e�]j�:�R>�u�'Z�X�]�n����7���O�B�����[�"|X9L5���_��[�I�\�$�xE�xT+�_'���'�W#�������ls�=S�I]���5�!@8�`�{�Z��l�u�ɆC�{��T^�%�P�b�����
��-?z�暵���y�i�����ô�ٿ��-� .�вm[�!=9�T��m�&����R����)�f*dGG~�t����[��� �"����Ŝ��y��	[�Eq);Eq?;��gw5v-��q��Ϋ�h'b`V�s4%,�X����:�^M��4�l�����x�?���`ad�vz71�+��[�j�9�ʮ�h��m���?t�qGq���;��}�� J��>¸�e9�xɝ*�[����
����{�I���K��S�S�AyfVl�"M��ګ��O����b�5}�z	٨��<%��Y�c9����+�(����k�"�Ec���������_?�d�NQ%)K���"��7�;��	}�p�o��s;Z�UM�]+���࿗�Z�J澒;z��j*<���"x����O�{���RNa��̞���b��@yȦ�h�˓@���E"����流�U��U�"�'�b�L����}G�y�]\�Qgwx˸���w!�/�����,[������3M���'�ܜ��˾��RC�yAE�]"S)�\��+P�C��/b*�j��H�FOA#�����Д��"��B�oJ�Q�˷�6J���|_�'������1ꂃ7κ�rW.5�#�j�D���:�d�~�򉣓J����
U��.7c]v�e��'�N)%�<�7��[���,N[e*�RU�S��Y��Vn`���|��?f�}�.k�O��m��:��P���~+��W>np$ϝ ��l��f1�1��?�ꬬRm{����hZ�[[EC���.L����˓��>Ś��
�QXz��C���?#��ݠ/��'�9���yg_���ƚ��\��B��ODp ��dҙI��9�z���R����J�S��x�8�H
 !N9����,Q!$����_�}�q������\x'ﾷ^��� ���Ϥrr�~Ӊ_ܫ������0c�}�\�˛K��o���3CKH�c��� �ao_$Z&���sx�ӨQ�R�yL�AB��n�"�k0-�&kB4�ҚH��dR!�R�n��t���t��g�W�*?��ϫ�0].�Ǡ^�3��Y7�D�8H�C+����H�����a�㬵�Ψ���#�����]i�I=3�?�Ou1k��_�B�qNl���3��>�	Zq�]A�ԉ ��X�����Iv���rD:|�N�[�����%�̑�p))c��s�%��f�w��}0�i�q��2K3Zq���cܰV>Ke��z�SA���~҈�X�A�A�@�Ќ'!U��8}~�Γm�+�qμ�%��a4%g�r`�w��$��n���|v�'�W��ii�(���0���l�%طd?Qϩ���X��w;��)G���u�� ���sK���d$䍴RB�m�2�as�'�7�s�-M��]��O�\&=���rw�re(IR��8G��k���Z�S@ �J�8���S�T���U�!�����i�)Z4L�I�s��v�f�˟R�ty}�?�eJ4d6TƂ��ؠP�p���$���8t��7�pb���]=/e�*'�oԾ������>�g���8� ��uY��墯�0ClcW+Y|�mݪ������+m�Yy�⭏�*:{��Ԡ�}��&d5�v��mѷP�Mû[	�B���x-�`R=r/b�`�Q�1�Ub��˖t���J�{-���F�皂O�Evn7���⌖���s���5vMi�|��|yM��K�s\<=O�Ѱ�O륈�)�ά�Bd�2��s_l���ᕋ�$h��^kj��W!�A<[���Ȳ��dP���(o��C�X)��N������*Z�O�s�GS�Vi�ubv������Ф��'Q���߼��x���a�ze��q�S(d��]����R�_)�T k��&@���M��������=Ro�{�z���TV ���e(��6fL�����z��e��,�[���il]]�`���ɐ����}����p��M��w�e�����噫Vw�wb�;�Ь��g�}�𞣫�fLu˿�	�� ��M
iW�ƢE��L�6�C�^��7���ӡt��o�0z�f���!޼gV|��L��e�ݳ������*��?�&�"� �S��Ǐ���K:=:�����:���Ǯ�b����e �,����2��1Q�[��&���7*�-�=ʗ��)(��ŕ+c}�~����w���y�υ#����)��3�᧗���f�k�,��"�Y��f�|��Zt���d����)�d_�N��j��!5�m�j���Iٌ<ts���5S2�s��ebK2�����_O(��)�Ҝ����_󞽴������B�^A���o>�$���I0�<�9eT�H�y��f2\$�e	$�)�EG��q��߾��5؎1������t����&�K`�v����4�P��P��ϳ�T�|�>	��G"O�i'�g~>x����o?|:��s--�����ز������K�"�Nt���<M�x�H����}w �ܐ��/z5ޫ3�;��C ��쑼��h�E���l�  Jj��:,��# �7<2���n?�}ap�/�V���Z���"Sj�{�֎2�܋�SE��UVGz7��bS���-�5���C���>_�a@�cE`�\v���qk���iC3�G��vu�P�Kq.�B6,T7�!dlZ2��[��3�C��ow�QjqV�N�J�O�K#
�P�8��~������ܜ��S�&\"k8���M�Eq���]��:-q�w5--����;-{t�%���vzRW��z׷�#?r���~�[��S�B��B� �����d�Qa=Zta���O+,n�<9���Y>�,)����|��ե�j� �螒�7����^�%���~b�2v���+�j���֪ݢ}d)$��!���0�.�Խ�.y�,��`\'��H�!�+/q�z3��X�m����4�қ���ƚ�����)W��ҳ���iɰ�5�����X�H��^��"e$59'Xk�d�N5��4���+��Nr��d�Smܐ*�� ݆�;2K��"��k|��A>���#?
�
P��j�6����/%�!�'��'�m
Wo�p;��"]���ŏ��-��+PS@K&�ޙ��U�XQ3����3�/�n�nG��eu'pLf_f��??ɧ���0h�0��p�^�$I�����������n7��`|:s|\Uo�"h-�J̱r��NLc����O˟�1L�w�2�Hk�$1�ǾüX��'@�~y��)��AD�b�!����u��*��Y~���&�N��@�����y�#z�@NV-+�2����ڼ]���/K��UR� �0��-u���9��ӛ�h��4v�@����M��t�l�?ӺL�@@pC��E�Ჳ���,�&Æh�S���[M��߱�j��2��톛`�������FhE/ː��a������k�k?b������] d�Cj����y�� ��H�n�,
�K?�IwH���<��'����^0r�,�=d���03a��U#cL% �O��Y�xJsg��
a]����a����Eo8��'���V����*3���B���J�m��4���k�x&0@�K9��	9_F�:K��I89��@6^�f�����!��ܲ�R�O��~��'mZ���^s�L��M�"&'�co�P���!"�s0&i�4�e?�#g�������X������O�>>G{�#���Y�k�λ���
�uha^[^S����욛�H���A|CpS�Z�un]�2�"S72��U���秧��N�ʊ%5���c��=�z�����a֭Xks6�]q��;`pmc~ӄM��W�k��<�h8U��@��@x��{�V ���C�sXX ��*�����I���U�!��$F	:�7_0Jz�NoP�<I��c�Z��e����T����D�C��I��\�o�������s �HB\X�UseI��17>!Hb��}�Q��f���N�<jr���{���h\x�	о#�uJ}a��{��~Bܲ3�������p)!�Y.�ڝt嗉V���w�ɘԺ�e��7߬�<��
N�s�� ��3�궰���U48�k�R6@����jp2V�����Q�q	���:��Ԅ��D�A{@G��6���%��yE/ry��f�j�Y"�[R��[^��f� \vݜ��ﾙ�:w����4��H�����I=���9V}'�]��t�{���z�����e�g����'dJ�s��ڌZ� ��i�du�4��c�U�^�iAM�7��8�q��9]m��		n�+S�7���*��t���	���[J���]�U2�͙��H�ԟ�=�%j��Ϫ�U��$�҉��p�ߋ��Rh%�d��^W٭p��j�c6�E��^���R��3P����j
��܈HB�u�`7���'��ŰL��尰�K-u����{+fgk]uj���j��n��NR^(ig����*&cW8���O=�5������nj��房\e�\�F>I'(ɧ|A��;8���U.TX�G�� �p��>�����E㴦����_�߫��C�v�&�e/dUx�� �&Ĉ������1�2��tU�*�rx�cX�84�1T.h�И��7Tr܉H���*}F��*O��AkD`��H��mv�� "��ma�7#�`JK\ȅ}�)�#�M�g8�wz��d��u����2�P#i��$?����'+����(�	� ��g5��rjt���![kC
j��OC��c"촹ٝ$0�GlJu�љ��@>������u�ʚ'��Q��Ac�L�=]�ZB.�����O�}�{��W.ke���9o�e���.�'B�bb�|�Z�ؽa�=�&�]��i �#i�Pi~�/Ք�3���"��z�85�Ҁ�$~�s���Lyㅵ�N-��D� �;: i�A��Q(ԧ1��rf����u<y�p~�v"+p�!��Y�i�wl�.��x�Y���Ǟ���*��8K����L����⠡�;OY��va*qb��x�.;�ЁQ���A�JXiYM�:���Y��﮿(�)���ě|�9��(}�W��6[w���]��Tj�n�<�\
E���VL��C�l�fDZ/�Q����<۞@2���Nȕ� ��y{�Ǆζ��I+�&�B^y��	����=�|��W��N�:�R��&^f�j!/����]2��Ef*F�nøl���_�z�с�kG���^æ���&�I��O,]��������f�j�`�� @L��L��`=����6�z�c�7���lk����w=������P��42/I|\�WX�&�r��J��=�'SknH��]�#�#��`5g�ZIo�U�������,�4n{��a$�x��U� D_���r�>�~�Y��$T������!S�wdx	�p���kU3�7���!M�\�g��X۵Ϥ�02�<��Rc�Kg��e*x��V�x��k��-æ��(lyv�@�חQ�'R�����d;�ɛ Z��O��V[(!K�C
~���"�2����ކ*�'��A��3U~~~��Ҡ�{w��?.�s�j�ڌ�O���ʞi�j˟�k�o����Pz�Y�%e��M��|�g�~�w��~�� '�| ������~
�EV�����..PS���)(���î��)��ޏ[ޠO��P�l��վ;:ظ��L�՜vv◔��.V��|�͇��:gQɆ�s��p��l��� #�;�o\Wҽ+*����RkZ��frh��]���^#,������࠽en�J��U�N�Wa��-���O�Qi����Y����R���(i��E��!�Y���)w���gl����.�X3ȩ���o+���3l;1k����y��=9/���Y�[������4fN�<����q�(4#&�׆9���[1��/u�?@l�2�n�a)-T��Ŷ�<nբ�����*/��)��Fȵư�8gT����_r�\_̉A^/j������4�M���d�_��{B�O��Dk4���mX!�#X��!-8=��z�Rov�_u~����'�L�b��u�*���'�����;,>�^��9s~N?�����G���PJ�q@�k���*k_�ytK�z��A���v���ѹ������<3���Ic��>������gv�M_!��I#B���!��Vy쮄�/���� <�cr����G�͞�=g@wv�J�G�$8C�!8^�կ�YZG�-i����%m �$¸�!�4��"wל@p��qL��c�4�2�C%�^���~��%S}iZ'�~�2���e�^�t�lj��Ѹ�E�ί#Ǻ�]���>݌;���˷g@� ��]i<��=z�\�Fe6�lD��ۤ�Oe��L�e̷ny�~��')���Y��T�\0|<	���f�H���:ӱ�<!������	C��a��[[2��ra�d�_�<TF��zhM/�ɚ�����GK
�>�j�(�Md�;��~�}I�އ�c��d-�^?]���œ
���p��0�M��w:JoF�I܁�a�� �'�j�&#��f���|��+��>�1y����4�TWk��B�H��d�- ������[��c=;��ޮ�q��r�L��L>n-���%-0�K��0F��3F��=(qa�%�����wy��ޛ�,y�S��7ȿ���y6��+�4g(j�ȅ�Ú�)!^/~���Bo.��z��#J��	���ʞQ��In��A��[C�\m��t�>Т�}k`ǣA�EF=L���U�=ј�WY��?0�T�K*AZr	��)�#o �M����gp�6v��v���(��Z���ߴ�1��o]R2����}R4q�RM�kh����<#c�k���a��e�͹�_/���팅���i����B��G���a �?��j��'� �!�W"�O՜��{��׳�u�E�pL����h�"��|��C�ū���s���=b�wT)�Q��`��E�y_�ʛb+��^�,�����������x�Q��Y*R٪�\u�P�5�Ƀ0#Uؚ5J�AF~�lf�]���}'���n��l�nM�?�tj�m��W�Z�kE�b��4����fůq¢b�X�{�C��E��"��_������<ҩ�l���]~�ۦN{U5!�\a{����5�]��O,�����&�X[!��U��bΠ���9Xk$s����2���s�?��_�aH�L�Vf_� ������R����:D�Q)0G�����s�����2�v���BI�����7���$w�� �FK��I�W�����W���u����+֞�^a��(�{w��?o���,x�w�	�i*��\	�.��]���t
֤����u����+к�|���XXřW��>/3%)qǖ���J[-e{��;�Q��%�/��0���Rg!���Xs"�n� �Fؚ����\Y�暰����Y�Fr��[o��X���m<Ɔ6dT����4���>y[ri7eiR���;�m6W�����-z�0	�%q������ ���:��O��,��r��Z����Ǽ��Pğ�\�u�P��5�3/�;?��D��B0�`���x�7k�1��&�[܇��b�]�uԧ�9�� �?���l����F�cOv1��~�s�k�eutһ�gMD{��������._�2�$v��l��ޥ��Ň��zȆ(#y���T�c8@X���n�a��׾�"q턮a�K���q���w��c����3֛[,��;e�J{��j�}s�+��쯐���)�\�?8���v�s�����Z�J��
�WwP��s³�O�G��|���_|�`��u�sL�bZ�R��l7[�7��᲍^�ƺqS����e�������#;�� ��`�훀��E�z��v��Q�qA��Pj�>ZFȜ��~BaQ�e��w,$�io=+��zE#�ha�\�k���:�NQ7pn�nnֿ�L�X�qQ<�m�;!��*�V�L;�*`4��u}i�MA]6�'�O�������K&=(ҵA:�� .��\�T���b�[
8���/�?J݌��v
�J�\.�#3ImD'�O{_���'X���)Rz�SO^J]��qi��U�^\�M`������7ٗc�!��Ơ�p�q/�]�%��(&w�A8���*U_���e�u�7oxp�<����i{ϟ����ַ3�uy}k�?>�r;�g�n��e�D�8�+GO�~<���DN�;G���g}��-�C�-�����K�5МO���t�^� �p#� ��'�+ɻ��v?�a�R1���|\�}E7od��ڜs��2���k_7W�<�Ț`=6�]�w���v~K^��ږ���^�0�����g��D����I{E�Kqý�ER�}�)Vu���*�2ހ����I2�Bw�/E���	���n��c������-�p���JV	g_�ٍ����P�( ���ԥzh}��>{{�a� о�k̨�(�g�-.�:���{V/�n���|���4=�|a1��e�˷�����2�|A���O�,HT�Ձ5Z�U�-4_	L�{2���B7o=m?ȇ5��1����/U�^�V~��u8��S�m]�=�zS�B}�߄1lK��j����f�p���y?k��Tl��������t���g~!`a���b�F-��.��hP� 6C-߈ƢY�o��=�U"�DU�,Rm�Ϫ�?^�m�K����?�{A;)'{H�x��F���)�.aa3��**��!�_��ˬ�n���^�k��
�j�p^������x�y��������rs�C�}�7�`iN� �v28��V @�1X\�Z��{l�bk�����m篣�����)��)5��(NEy��+�Q�|��SW��by��!��PS?fR���K����)j�@�]!~C��c��j`������a���<�%�6m3��*�,��P��lN�_⊒����)F2�t�� e�1xE�-6��"��gա�O��!/H��B63ǍΦ;�#�U���XJ^T\�(:��k�w�iM)Ѳ#ϡV��O�nY8��]8��w�H|�v�T&IhYn��y�����>�]%�FEԦ`�������B�J!�I�nW��0��k,
��>�b�W��4媉����[(N�ӕޠC�iсs�܍IS71�-rḤ�-�cg6�uܵF��E;g�FO���n]r��Pi��J�����!p"�pB{�v'櫫�b�>ʭ��˹a�K�Q�4tu8,n�E�6i�I��i�R�\�}Dy[X�(9K�ӳgF��ijD�f�,��b_1�=��X%�F�tu�7Y����ެ�/����=���;���&38],n�ja��/GC�!M����}����U0��L2=)j<�s���l@����Ίn8��]cYą*}�p�x"�]H�<<��c����| r�{�H�����u�~�ǾZ���o����'�ko����t��"�T�6b�,2�n�Q%���yY��[����A�(%�R��v��$h]P�J�ۢݺ��ym\v̈�F�j�qjH��>�azR�z�޻H!ŵ����n��Af��5����c�렛���g���g+nVg�=��z�ُ�h<�}��o�ie��R�S�ɯ��֚c�Ӧz1����O
�*,>��F�K���u��b�s�\i�������8FK8ED�oyڲ�)�{eoɯ�X��8�o��<����;��_T.rO�7��]��HU���??j�����B�J}}�����������JPt�����������O�n�.}o�x�d����Xþ� ��ӡ�"��$*�5�h&�,I{Ķ�E����Z������s���~9�O�b�أ�5p�w�<��e�W�#sW4���R��u|�e���]�>wZ�!~��l+vJ��$����\y���S�]�=�%>��}=3�����CW��\��M��ؐ��.��p�l�z{� a�H�s�Π��[}��+��[�$�]��֗i���r��8ĩK�W���u=tZ�o� ���N��`Ι�4��<�fH��]�~����p?�vP'|#�X��y+��{�e����}�9QVW��~S�
���qlz	zj\��9[_� 9�~��	w��)'��=ۙ񩶨>��r7w��:9����	�7&�i$uv� (��&�N$��g��˴E�%n"���&
���(��ؖ�%TE����'�e�{ �|���y�����\�I^&���55��H�y�w����Q=���Nn�o9�ȐL�R��iJ��Ô+�-�N���Rt�a�vc�aWY?Se(K��b[��S�#��{�c�R��~�>"�ya��Ɛcr��M�NՋ?�%�_�h�j:��1z8�9R�������]�6��aI.ʣ-]r��D�F�G?�r�i,?�?����p~�DٿN�J|�'7�.F�o��T�G�ܳc��h�NZ��}k�jƲ��^�����i9��(�
��Rby��cQ� ���9�0��f��%�m<yﷆD�D|�Rf�W1��������C�-�'9Ba�����*�eG	��fmuC����E����WC�W?Ζ���������eҞ�_!5*�mnY����|b�s>�i�ׇϋ�$Oû)�[b*a��5�l��1Z��/M�7�=�1�[if�1?� �?�@�������3���U�Q�e{/�)^~���!ɬ�<�A�������/e	�$�k`�SV�)����x��d�㽸�v��?�}1[`�� ��V{sHɥa,3��7�쟧�Y�$�te��&��Z��Y��5��'
>F�L3�-K�{$"��h�N}��0�b'U1�\�
��[�X,<�����X��L--�x�j/Q�bˬ��44a~9#b�W�o����6������j#��:�}�답>��S�!�z��rߪC�����;g��J??Ʈ����]��}��O��2(3,7}u��b�[��J�E��=���Ɉ;���������������"HI��HHJH�4(=R�9� %��%-]�=� ��=CH����Ũ������ٵ��������㉉��`̚CC]���ނ)��>Ԭ��+��u�nm
�z�T��ώ+�98!G�7墼��D�Wu�P�ZI,b�}�ܜB�G�"P*ƛ[khՖ#�9A�i�w�W�~@�N1��/�f���v��T~�D\�W��%�	�t���\�>�ֳ�E��K����0��>�M:�]r�W��9��
��7O�w���֬�%D�:�"4�곏-��uW�d:���+�B��;�Ҟa�P���%;�L�PÄG�%;i2��;B�YZ�S�0�����S9�	���{Duy�g�F����v�'x�Ǒl��[�U�h�ƈJc��^�l����x����B�sб�>��͓���K�jW����Bi�	6`3{����<m����i����1�-��S.R�NU=B��J�b���
,�Km��-H���z�ڼ�N��eG�Oi�N��I>)�����b���\����WM34�Ս�����s���y�x������������QT0S(q�\�S�fZG�P��`ڽ��S��F_/�[����y~��L�����*�|�>k��;5�`����-���?���+�Nʗ9$K��0�Ҽ���|��I�l�qR�1�a2r�*\V���8�8G1꺄�χ��!D�󪿊�˕�&���_5?w$HYy����A���`�u��jN�Y8#P��iX7稷ҕ"ܬ!�H{C��$&,���#�z��:ؚ����<�slrSxF��_�ݒ�[R8�I>ۈ�X˂���w&�����<7�o)`!�\n�����tu�VW9k�I+7��f
E���½��h����Taާ��n�	����	�Vׄ�䧻�F�=1ױ3��b�ڵY[g��J�����O>����?>���LlN�	�)�� ��p�]��i�ZV뒏� ��t�ca!)��\K%$TW���S'��������	��
�Ɣ�?Ot��6|:ퟍ�k��x8���Y�]Q�����w=1�����[��&`r�/��ꇓ�%��O0�ף"kK[�ԉ?j<VU^gꔶ�?�tB�A
�k�h�v�v�H߯�p9N�P6��YH�H��*����.�4(��������z�j��_C��Ǟ��px�q��J����l��
h#��I��<�(�*�k}���1P_���?P�u��ؚ)�@�2&���(���D�e�;��7R�Tb*��v;ڳn=��{2���p&�۾\�uՅ��/��E�1���-��[z���lI�x ����f!��s�b\?��]D�v%�2�{Y��3?��M�C�7hw��B��(E\��YMmJT�f�����j�g[�� �-c�=�@�}oɲ����ؒ���7K�m���TЯr���_�)���'7y�`�1�{_n!�b.7������v�N��곣=����L)�]��]e�j�[y q=�ӓ�S}�͘/N���ߪN�Y-��ۑ�&5]�Z��'�`�R����%m!�u�Dh��_2�5P*:,���7�QE-$Ϲ
�%���L���6<m�Gi��+H�̶}��8E�؂����ֳ�x��� �2\��-݆-T�P�^�Ic���~�ypa�ĿJp����V��l��Z��*��x[o�G��L�m�nt�����`<�D����9w�|WУ��ä��R/(�p��@��	�2��q�䇒��|�U@ܟ��l�LԄ���iQO?��w��D��6nX޾�?��m�K��XK��B
�T�&�F����b�2���*�������֋���
�CF?�ص��y��G�E���.�+�p�jm7�<�9�;\��ºrԿB�uWt��\H���ٲ�!��p���,��dH߆���UGxK���uWQr�n�(R��o�����`����k`z�:Yz��MTG��j�6yK�\��v�=�a�)��٦]���%3!^�p��!��nJ���<������,~�4��y��.�LyN?W�r�����<���-�@u)�\Ä=�Ҍbǉ3��+��
SK0H��������7�BZ.��f��q�9ga}`����S�+� �SG�[��
:\���}����X?��/o$� xT��s¨�M)����q͍!��$=��}0��;X��.�ٔ"M��� ż����(y@{���y�雚^�{������?�v7 �Sa0;ah������N��+5A|��Q==����[��� �����u�.ɂ��x?�eW�I����0�H���@������z��j�k�[��U9	S��ò�v����ʼ!���G��V⨧RS4���ܚ��� 7Յ�����H���>l-ƈ� �DLJ�3C��ٹ�Y
��Xͼ��͖B��,4����,�IXj�e��lx�ѸV8#�p�0�Hd��OE*�L���2�Tv�ӂ��P �wW�F	`�6n�PB�=,dN��Ԩ6�ߕ;��T0\|���}�%r�Bh�E����N�Zc��L��<���*��k҄��J���E��L��A�X��G�z�Dl-������n�v/�3�����¿���5�BL2x��?@0�l9C�C��C�ء�t�kQ����)L)�����[���'?P�@=��˝uq�w��x#��5z{6uua5�7ר�h�"Q�;ekql!	&ۮ�1���ڇ�U�6
��͓�(�/�r������|1�
�T�R&h*�Go"{�-�.��!m�*��q��e�9s������;������X��ؓ���nt��9�3v�{طg_����O��eAuk
)ɋ���>J+/v���:Iˑ�����i!1/;ZH�[�=&�&z"��^$����>!|kF�J`Y�R_UQ����r�ϲ��/#Nk�5��i_�9�J�(�z:�m��'0�с��m`�x �[��輾�UA���F�����X�h�:{�RSw��H�����p�g��{�'���_��p&J������O6t�|T�Dp�ڼЩ�os��3�s�0�<!�BEo�BtS���>�T�蕟T0�j��`���뾠{z����H��BxeL*`T�✥ɤD�}�Co���`�>3�cgH7#
�>2;�����+aU}M�ߜ��(����ඪ�$!��z#r�d�4�)͒��S�f�=�ϐS�<7�[?�1<
d��B��'��G_���C�>�U���.����h�X?Q��X���7�s6�k�K�#m��� �����Ǣ�]?�g������R,7K�}�T� ���3g�_�`�<�����A6�����(�3Ϋ�W�nx)������!;ȸL8�P�g����{#��6᪳�[�+���ϭ�ׅ�'��J,'�������<l�Z���oj0�	jĚ���ۋ�o��R%jgA��z�R&�ٌ�ύ~���5�Ï�a��<�Px����:���JOBv��)����۳�RK�����o$[zj?��'럱vD'+�� ��r�� VC��C5�s�k�*\��0��1hгhG� ĩs,	{}���#�;8s�١�� ��a�%�9�Z��Q���=��%��B� �?+h�	�
�[��׎aG~�2�j�aM/LÛa��N��v�;�'ά\�����6��ϳw6=~*)�[��T�>���՗N����YT!\����NmSyUխ�? ���+�rt8�^oh��8��2����ӕ=m���-�1��]AM����Z�V�_�^�9���7�h�l��<O?�{�s��R7��܀L'y_�=ш[��I��i1�}�c�|o��w�Sq�T���t��k%�.�f�@/��8��<-	S�b[�-�O.����%Q{�]�r\�W���u{�u�g����ȿ֎�Vo��>ٜ����.{}!�˷#�-SͷS1�#f�������TI�D�O\�0ơ!w�W��ok���DG�=9�3��9rF_�~�_WB���x�M��Yo������iY�\#�������?���n�+x(kD�����)�L���K^�B����S}�v;�&��/�H�I�u��e�:7̷�l�AαP~��=�f�؟ӵ/�޸������:[~�^;h}f�9^��(�ɹ���K�?�#ʨyN��:Ɯ2?%N��yo7Ґ�[޸K&r!��'���U��X����[�ԱY`��W^�?^z��DP�9��?�O�K�>Omðj���#�\�hQH�����9A�Ycn�?6�5�~ZKfDu����A�'�?�lqhPR�?�\��9�!ar��/�7�#���B֦��b��A�X�+w5�T~[/��?U
,���@�Q(<��_<3��Y����v����~w�O�2�f�>�tWE?;�r��Y��m-\�\�ԔAG�������+������&���[�^Z�O��d�4�77*�E�^��'Xl=�/7TqS�G��t�N=L�i��ҏ�ԗ��?����&���k&� �������$����R��cg����[3��]�d?z�	�0�)�Q�L���xΠmZ�l��>"����
�	 �y�5Rn�e
�a*M����� R�̢�~�nE�h��']�`��2�U�q]ڮ�Ʉ�J�YN8�K��~0��r����"&�]H����s:^:�JМ{�����5�	�f_�(�ďo�١��{ہ��"G�~O�B���`��(5O<�w�t�	���Cl�Ñbs#�~CB
\3i�'����:�ݎ�t���Sc3-��y���x��z��Z�p�������׽b�4�qR;��R��G�ʪk�+`�i���xCÂ�}������Q�Pr��Q����8��oU%T:��wF��X���R��:���WR�`CF���-@��Ԗķ�oL ��LB��`�)�:-YY`�V"�l4�g��!w&"��(7���UJ�J%ӹ�3S��-��b����g����XWL��7���0k@?�V�M�0SЁ����i�N�������q�2��(G'J瞕n$nx�@a�"�@�'�^�opT�
�g[w�A֭3��n�,���l*P)��-d�:]P}濯6I����#���M�(�����+P�x@m�T�y�s$'%�	_-�>�T����r̢A%�j+�kˁ�����ّG��zN�O��P��N"!
�u�[���Jv����Z0ۤ?�������N� �����{+�w��&�h�M�o��^��W:����~}��I�soyU��ң1RRM�;噲�ˉ��x�%&v@����UYK�}��-6����{KD��^�D5M�:�`���i�p^����8���'w�q}7��.��E�[s�:��v��̭��=�v���lC�nu���>��;�_J�^~Wox� �L���kI\�4'�o��q�F�o(�=\k�|#�s�k�D��̙��s�;Up�Ǳ'��5H��'��H�d%�D�u�i����hJI�> ﬃ��?��Xn<׳�L0�E�s�쮤u�u�Ԏ����E�t�[��8�8o�v��:	�NAĤ|ڧ �Q�f>l���x������Y{=��u��b��qI�(��m�Bph0�@�st�g �G,����6Ur�G����ߝԏ�w�/��a��p�_�H>��Q����B�
�{����zg�7�@���e�:�.M�L|K�r��g'+Dt��T���=�ε[�����v�a��\y}Z)�A�2G�2[��v�~bΝ��-��Dv0uL%���[2�� �]7bJ�DJ�vm3�2z�^�OnΔ��D3�o�ك���!k�����K��"�+u���F�Ƣ��'����B�|���{i�o�����J	q���w-�^�o��F�|~8��Y�����������6��k(�&��d�~, [�P��?đ�-�Yք�����-L�C�:z`��pɟ�ʛ�q����T�]'a\�j�~�����T�n���௤I�yOsi���Z��΄��#?Blсd/+d��D�K,$�f|O���Y��% �����+m�B>p����o\:
P9O҆���H�����R�~Ş�N�O�(a�y:<����!���䵐�;��R�?q�t���v�<�+A�`����X���rH<�A��-��DI��^����{"���U����_?�y�oj�߂ol�f���Be�������c�Ё�s��T�I��i��A)mǽ�������������*���Z�zL�-����:�e?6��q��QvL������=5�^��i��@ӹ�Q(�u�5��|��u��
ϻ)e�ĥ%�th~r߯ukI@I�鍧��>��a�����3`�{oG�q�B�J�qI_#�������bf���l�\�۝2�ӧV�Å{^o�hI�hˈ^a`��G{�oAv~`���4�������Tk�O��d*h�ϥ��-ޭ�A�Χ���x���t�Y�=�%K̯��0!���eD{[����h>ˍ�yw���ѼKD^��Ŭ�]�Y��Y�<���t��b�[MR+�#L6�Z�槩������i�j�A�I�1��e�Z�'������[���V~������������S'���<H-9����>��ʈ�:����e��j�W@L���\��w��7�8:2�]3�|y����������Vt��6�pI�u�am�J����HO;��d�<�,#���{"�[�u�܇��:�\�z����;.�g��pbr��`Ծ�Q��h1��p�#m�|�~�ކx�:�75Z�1����+��vkb��p3���D5d�;�����=��]�/vͯ6v"�3���?�����m�e ��@�W��鈍�5.u�=����LΒ�p,���d�<�7���M�t)m���S��=�MŹ����f��Ƅ4Ӕ���	`+�/�n�t�
�`�;�*f���J<U�nz���i�'���X�֩x�s�^��]�����������b�~׵��nl��CJ��7���I�o������"�,��XO�m�Z���ˆ��(�O�[�*�V�Hm��$	&�)bw§^H~��oX��{G�b^�a��}i :`�e���H�x�����]�)���b�;�P���>���������ӮbSپjލ�4U��Ԓ�j���ai�̾81ID3M��~�l�f�R�M
:��3�b��rxO4oC�~pZ7ϝ�}g��.���2�+.�1�j"�s%/��dp��6��sm(k�!�'�/��`!��L7�a$k�R7ѝ�=?��}-xj���w�~"�W��l��ݴ�tZ��@�4�f��Gx~�a����EM���uh�n{9�(��<"�N��]��^{q;^��sf!aё�q��W���?�������&��e���H@ ؠm~���F�K�V��`�4Y�Dy�'q�\C�BU��S�̬~�%�'�:�X����Ǽ��f��9�$�l��_���g�J}н�{��*Y;���"঒�͌%t�jP��ܽ�9()�r�^��]���o���)�L<S
�V�óﮅw�W�gͨ���C�O��=�isf�݂.S��tzl��p�<r&��t[��a	,�-7D}8��'.�)����A<S��9�V��5�?>)�e�o�z�zj��@��\8VQ�V"�or	��E�7�{�[�A��l�*~+�^�+Jz��j}����QǴ�e��uR�Ƚ���
̈́"����<Mobvo*��±�堄��n�[�l>��Z]�<a"&{S�2�zk3VcFc"?��=[k�Vҥ7�}|����Hr��0z�B�B���s��vȏ�>%>�bכ�2�u(yli�&�ŧ���]��Ah��$M�&�`V�c��W�{+���2oޒ*��ϔ>�w�m��U32e�>���c�<��9� Dw�S(�#r�����ܵW99*�B�-��� ��VT����M� r��m||)�1��oϨ�)6�ų�6#��nyƪ��n���x���<c� }���+��C�&�r��1�k�	>�G��j�Rl�M��6PΝ��P]Hŏ,���t /���0huDq�<���T1pf�1��!���k�����'�nz�Ar2/�^z��X{@t�.6��OD���򴗎fo�
�B��+��o��|?>�d�Mu��8B /�`[/T��Zx�~fH�W��c]�'�aq͚��س��J�%B,�/�
󋮏m]N����-�9�^! /^I0�A�%T�IV\ a����\\�x>�trO��V|rd5�����>��:��#v��؍�4Li���ꋦ��B���]s��p]݆������7����K�&M ��$�)�:�ֲݩ����+�� �A��ow��S0��:���ra6k8M���ˏ��⧹YK<d�ŏ���p3��	Z�����t�i����'G���!16Ec/�����8�i�3��O��K}��0scz���j�-�g���c���I�Y�}�����q���5Ua���V.��Uu<y��.��Ժ%tg���_��ޱZ����K;�G.v�z�8gc���%LI\DԷiE��N����\~1i�D�����͖§_��"�'��0kY�ʗ��E[��a��
��|�{�D@^#'�&;"H^-ֿ�p�F���I*t9R0�u�=+V� B0�ɋ�^A~@u�F_P��,���ZW�\G�`�,RJ�T&���R��3���aL.-��x��[_���u�!��k�F����K�	G����/_�a!��vśY�bc��9%�p��	�;���j�k�%�~.���J��ǔbV��	1����g?�Qk�r{]�1;zd+w �泑Oo�܉��G�O����:��=ҋg,3H�+�[4ٞ���B$K��Q�F\��o�k��7�E2_+��w^3o8�e/���f�&�P�6S�.H��XMu��nt��z�������vw=��ͤҗ[;��vV�r�խ�j=y��j���'���c7��L�᷅ܺ{k��A��P�9�z�@�?5���q���Y���a����_��,��{����~F)V/;*���8%��lx'����w!����Dt~"��5���Z��殏vs�-�����q틍�Y�X��[�c9�b�f"���
��@��-W���[k����c^��E�[9��F�
:FEE5�ݸ�?O!Y�}���g=�g�����Y���m�vR���t蒡�=>�s�WͶ�ysF��;n[��r��F]ë��+ncF2�X��U��*������'�+b������Se�9 T,��c�Zߒ}��
!�}}9�nFJ�\_x6����o��\�m�o���Ǯʋ�dep�3�˩V�#.�����䟒%�W٪4��k�B=a��|/xX�8���`��o��)Q�.��t4���{Z�i074ѡ�o�6W.�'�XG��S�*t׽Vg5�"���s�Ǖ�Է0ou3�~�;go�Z�
�'�c)���rs@�+�'�������E�x2�m�	����`[�p����@M[,���N�]}�k<�\��c6�q8Y�~��Zo4��O�e�a��V��h�ԡ�U��)q�=�n��O��x*��w��k�L�7^�)%�|�d�g��o�u~�g���HR7����"+�	M��>��R:f�x��RK��44zEV1jg��&�w�t�^W�ӈ]lZN�5� &e��Fc
�#D���G�%���ORDr�W1-D=���ź�.*�)l)Q�����/�,�V.���|�ǩE<����J�~�|�v�ԭ����;;�"ts���롟���{�����`u޵��1��>1^{���t��e����5y�v���G鈆ww�v+�AWe���O��b����ۃ��|.:¨��3��U ���78Xߙ�-�:�KW��M�4>Ӷ���ܟ�f���Q�J���F��'��mv���6�i�S�23��3��'���%���v\��ʈl��q�Jloo���{�"|j��z�%�~�(*S�"뾕��{�+�2��iz}E+��Lt����X����p/xΒ���ՙ}��(��j��-K U̷wL����l�NX���b��U������%�y�'�,V�=	�%�9WQT��v@aog}�R�����섰)�<���� �v��H�Z9�=���ɬ�*Vҫ�丝�O���\�nE�MG�bx+D�oM�������eS$����$^�]�{^iVF���-�?I��%<�J�h�YY�,�5+�./�n��F�z�q �&��Ζ$������=T]���e��e7�{�Ǟl�6��}�Dn6����iz�GR۸�'Sk�s��k�������7(hO	ҹ�S��GS�`X�Ú��Z���-'��`�_���!B���0CB�=cR &m==����~L[��|�)�> �����g��Dm�,j�8�JU��IG�Uq�U����=B�K��U_Hq �P��8D*��&7)���]��H{�X� ��xTHQ�a���;h�+���h�Y��+�����wA���A~/��rߖ؎�GHQ+ҿ8*R�m�?U9WI�ۍ	|���!6[99��iǷ�5+Z�f�#��w��Q�o+������V��P���^��b���[W�7_8K�8����/9��g�qO�����8W��ۓ���|B_9�|������p��ٜJ�H����=sxO=��N��t_��F�Ɛf#��˛���F2mw���o��к�6K׼�
�f�&;e��p�g�ՙ~E��FIZA!ף��������r=��d%ɿ�R���љ��	�lh���l�ڷߖi����KA�.��_Y�x����W���������%CہgB쭨2�/�H�B��E�6_�u����Tb`���(`v���뮍�z���"��L��	Y��/��W[]�6�V�j�+a�W31c�uv|��:&�=�sMl�� ��Q �;+�m��)U:ŕ�2�\n^<E����f�MS�ӟ=�mc�$�Ӗ�ČI=
�`:�@������a�U�$��\V����ǉҹb�K��d��=ϧ��j�����Ɯ�%.�ŕ�ǐ����q�V�Q�4��`wȑ��6��;���\&=Y�S�-~3��@�^?4=���iZ�.jx(V1��4�)�0�&%���D)�}ەC/���:o��f��d%�r�B�0��1�>�~��y�t�*��Z\v��DEM�=��g�jĉ"�YôB|�X�3M��4���Q����=R1�e�zMY�������B�y�_�-�d�����3����g�����=tS�ڍ-�E/9o� ���J�;09oƩo�^�+�l��v�D���`(?��8��p�i����&Ps�+ۭ���HP�-$¼�W@���ћ�1?��|G<���Z�Z�b�O2�(�bV6���|ixnA�����+�s;�.7~���O>�-�d��MJ�'�_�be��NwY>��uNuR�Wy��Ui�?�@{M.z ��$�jyk*����ے���1)�_F�If�s,���	AFo���U�ʤ9J�ȉ�E-�a��j,=ėZf���V�T`nA����l�L�O�D�-�D�Si�c���n�#`x%�W���Ԉ�]�$�Y@�z%��Q;c��r��5�t��#z=���Ʃ �����Cl��o['�Ὣӻ]��
b�YaݤZ�Ӣ���O���E*w��$�W�ަ�k"���������U����p���\�d�	��%���D1�����C��Vh}���|�;P�5}P��(3�&�9ޕ5�s:_.vqq@%��ݟ�D=�WLsA6�vYF�F�S�lO)p�Ǭ��%���$g8[\��%l�]s���R�7�E*��ش7����1_�R��_Sbu �2�	����=̕�V5��::Sl��y�S����3�[��%V	�ٛ�$+��{a���<��g��j���|>���f�?��sΚ����i� Q{�N��bO��52����Y�8��4����N�l�.p��D�%vc�������@��'�C|�><� �`ܠSc��"�M)E��m| ����Ø��̫����,U�9e�&�c��a����Cb���,�C���\���œg�E*�:�u�Iu[�?(L=V�x	�r���}��j�z�ԕ+F\KmAH ��sN����f��Br&���[�yA�/��,P�#�s)WF��G��s@MO,�;���H���d�^+���,�c$=��V)�r���y����iI�0��X|xU�G�8p��˕WJ�:��][6�&�q�[��
�.�1�7q��ӓ��3���W��<��0��S9��^��&}���׹�Z���b?�kx����5j��N�:���Ӧt�N��ʜ��Ҽ/#pi=~~�<����_�K�I�ˏ�J���3�?8徧��8L���:��O#p��{��kٓP�ƙ2�Q߄{��=Oݧ�#,i7|�3������{�Ov+Ԩ���+y؂���9�1���
�e-5�hM�#����O��O�paJ`))�^�<�K;Z߈A�HI��� �ۻ����ݒ�"�n�~	��oҬW�.1���Mή�ۚ���0�٪%#����Bȷ�nǊ|��l���_��|�K^3i��u�`����h�mد���͡������	�� y���Tr�+l�s��I�ҹ���Ԕn0��72#w��c�:r��YI�t�.xV�u������:���)�$������fJ_B{Syzr�ZO�_?{x���j�lGCC�2�;虧��ӏ]���_��|7e�ڢ_S%#���������e��.�wPL\ERr�UN ��+Nz6��I$�-5J
��������\F�,��R\��|B�R'\eL��S����u+4�t�&q���mӄ�CS��0�pr�pA�aw��B<*�5�;1Sͱ����?��8����������٫0��Oޭ���k^~�� �D������U�2�t�ȧ2h���V��{Uy�oʥ\�a�߯�|��A$�/G���pZ��T�T��G��jѢVW��Rfs3��p���}�KE�6�"$�e�i�d~����K\�&+U����Y���{jQ�F8���ื��K�mq�@X�˼]��Y� ����#!����D_�����/�+�xl&KKG��q�E�wZ>��xi�-h�j�9����)t����P���"}�gႷ9�l�'�i/�vJ�U=�đ�K���]��r65�$&Yt$4d*�_�0,ZM㵿�yd�>ttI�NI�Ow�css��,��^��]s��B_s��^��J?�^z�.F�_���d5�Y�4ltm�6�(�yd�:6=)�PI��}{�2������	�c���eR�]����nk����Ϧ~�k�Uk3�������䱲�i�u�G�7.,�/�_���j!�hm;��^"�Ewz�"8���
����}�5(���8��޹3���{y0�Fd�M���������P���j�	�bv�P�ѕ�r��������e� ^š�w`�]h͒��d��e�@��y!�U����d����v$qGy�Y�V�{�y�r�H���. 	pE|44x�\�,$��TR=��\i*l2%|�pI���7O@���0%��i��/�M��xl��?ߐ�+��	�F��HI��)���� �Z��c����M���D�
���ߨR�ڨ���E�/��K|�X����_m��$�FI"��ŕ<A>��}=W�$�b�����s�yhx��|����$^�TЀ3�G��_C'LUk�]NOEWVJ&�*�ϝ�G�f�qK	�UXx��&⤰q|>�7� t�X�� /�	K��'(�Ջ �'�����0 fE���^���U2Q�d�p��H����,�^OZO��~x6��(�8����M�y���|��!�M�7l����(���k��|�H��瓩���	��������|+z<��i1��Fr�P����z{ŕ����⋟%��;����dF���q��uqq	�l��^�i���/�W����?"�X����rT���dTAT���P��l6�Qq��@N{ZQ\�`��^�������*7 ����%.]��4��j0���?s�?��+9�;�_��ܘ�F�V�CuaMU�� �:T��o�G����5�[��_�[���m�����>Fq����d�w}����1ߩ��s�n�߈;1��T�v[8=I��j�������P�",۵<6��$��ĳ��	l��$�������z6��4��.���}��(��#�?� ]Q끕��b	aہ�Y*e����5����ȷw�D��:[�L(<W�sw�Y�&�I0�� ���#5���{9��C20���E��.Yj�|��?4$�8�A�z����_��'�pm��1_�����M:_*
>.^S�Ӭ�B|�-��4<_�fQ�kIn�_ux�8u4s\
��g��.�5fA����з�[�������ġKU���
�9���t�[�.�+����w^Y������d@<#�K��*K���-W0��܉��}~Py�zN��o=��#Ј4A% ���)���ܦ��.�����O��چ�*
����c=@7@�ݦSX�Ov�t3����4Օ.�m������)�uG�f��/�ʂ < ��()E����j��P`�.�ufƹ��k�i�Ai+%��t�
���>ʛ�����M��y��8��e=��Q=�#u�x 3�
���h�r�R~��<C�!}g0�*��mv�o4kT���ʝ�٣�8����)+H]��پ�ϙ�խ�!� a��8�����M��l�a�P�^�e�`ߝ���������Ĉ}Tdo�Rƣ��,Ϟ-�rƐ�>5����^��W��嚴�����tݽ�=��A;A[z�5:N�{ �G|~~8����|lm�I,_�n�|���U[��B	�����faSH_W�W@�1Dș�;�l�OlE �xW��Y��ݒ���y!��r�o�����E��]�؁�[�|���z[p�M!���=l6}�q�%�{v��}�Q�S�[� ��<�E'g�x�:�v��WΒ��V��\�EP��յ����Q�~2PۥC�j���<YnN;��I�0}��ꖼ�� oB�Z�E��P��%����:.q9���S;<�1��3�x#�(k�&k�yB�vg?�z?�Ȣ~��ݗ	/8n�o2�c.��=��XF��c���T/�+?�E�f�������}��J%X���<P[!�x_�4���O���R&F���_K�C����6ɶC膎���վ��ڙG�߫�/W�)��ssm����3M���cD��Mx�ᆾ��x�ߧY�6�����w�(3��P�z"%��&�=n}߉֦�����^&H�8s��W �gΟ�ן����d��Z��;<D��6~�핇r�ۜ������بv��aSڦ�v5��6L�Cw@� ^�� AS�L�	���H2�9�0�a��_����]��T#�a:��!K>�8}z�ɻ���W�TuO��By(	���=�����0��B=̐y�)G{u?	����ke�Ҕ��Q��-�S�G��h���|�)�ph����8���O���5�.�� Q���i�'F��*mD_%.̺t6H:��h58uE��2U��F�|Bdn�T��ƙ+�nw�A���%WW�)^'ә�� "8 ��N��G�:��8�{Lu�������^���0��L%�OIt��� �L��s���	��n�?qF3�{ߕ��b��
�i<;�j�^�]��>�O��I3�~�XF��'T��re� ���5߇Osz����M�`��5���ڼM��:\*��j,.D _�q�K����Vpa#����Ҿ�`�7�t�?��.�$H��cf��=
�S~Y�U�/}rc�L=?4����y�Ϻ�.h������C�Sڗ�0�j����1� ��t �w���87�3���՝$]@��||
̼����=�H��I/��Pxz��yC��{�^Aݦ�2��_C*H��	���z��{ۻb�~����Z4T�a�t4�3��:~X��[�Q�QUS-!4����N�eX�^�4�~Ėv7a�z�HC�]�
��i�E��O� ��,��{���0��?�H�<Ld�i�fFH�ȳ���#+R	�w4�h��prds��6>�����h�@�
�����tDt��(�wPTÅrlo&��%G�dM�e�b{���̻�7���C�us4���a'�Ya�	͵|�G�Z�y+���b��ɶ��]�7o��ϑE��Y[Uy���k���$�o����y�0������Bl죔��>>�_A�&�ʺ�6s�V�~M
}t�nA�|·4�9i1Ub4�⼢�q�����9�ǖ]_�ϩ�f�w��T����y�@�uE�	YGg�!�(����'�ä;7���)�S�5$P�i =�Sa�.N=[�cd��~ ou�<{��n�4u})!i�1ȱ��v}k�� �ӭ"�t}��D�ID���2����Q��O�w�G��W�'.Z9��j`���-�Ç{��^���n� ծ��T��s�����/�4J ���`1����~�Y��as#�(�HMpE�Uy@�9�w�,��L�aep��~��y�!)��ʬ@��ڸS����e�����f���D�X:h��N��0��[^�?�m8`��OdZ�ȵ��a�˽�&���T���eEo.z�e������~���\t{&��I?{,�ⶩm?S��a��p�{�m�V���OB*"~\ Va;�Z��+��D��D)��Hn|�b��F��b�����k��d�8[�N,|<���<�` !�[=pۜ�е]S�pQ)3���-��@Sn��9���X���pxo�z�6P˶.����]��u���%\QԤj��͚�Z7����y�b�	���A�q8�t:�)\gum�9���miQܦf��w[O�E>z��L��x����X��,�&�|Ą��� �E A��߻UU[��S��eEn!�)0%��#5EC:��"�nVl����<uM��kk��3|gxaJ��rF�C*HL\kg��m�%�3iL�fI��IG�r�/�M� �������u������7��o��[M$�������/�V��В�o%jx�g{���PQu��0* ��#��%"�!-CIw�H��t��R�]�0�4�{�����k�r�b\w�����>�M��>a��\�����;4z������q���Af����kWG2��/��&q@���U���s� R��r��i�u}�g�(�,x`��HL5n����ʿz$��|
ra�mW��k�i���Uy����{�U�<
�a�^���MVFB�':��/99�m��=��',��,;˝����t[��wB�]�~!>�� j�jj��M�a^,��/�%������\�Ke������6�$�E	B�Kh)�z0��Vіc曤`�lޣ�X7D�Rz�qӾzJh�8�4�7������'x�������Ez��%��q�p�Ƃs���a�-����Ы�r��ė��004����7�{*���U�A���j����^{�#��oU��	S��g�����|}��s�KI`��� {򇊏�l73�yF2O�ZD�Nd	���VA���5����i"<±V��9�f�4�d���J�vm.$����g��C�`��on�E�^����dh�*��n=��If�I���j�B�gw
%0�l��E��3��`6��J��^ߜ����b5��6��[P����"��D�p��h�r��ʇ.��D�O�5�4���l2ūBz��Πw Aۗpe���5�Q>,M�I  � =T��4��\.�Sܱ����V���<�0���q*%���W�� �����-B)(�;ކ	���u!�y�
j�w>�L�1B��v7m�h�y��j�;��:�V��Z 5*��KQ��j��Mb��x�՛��G�ah�S�9g��k�.�?���t�H�'4pp��(��&��Uks�3���͂�n���畗	8��w��]���r}`���K�Q�n�a;	��c�Y� ����w��u�����uƎ���8��7��z޻��_��I�Tu�/��qWO?��A���z��ɲ�u�^yv�]aB�3�:���;�ϙz}�qx�������'|;c	��;o�������/�k������\��=���Qz��G'-T�����}����Uߐ��|�U��l���S�0�ǥ<V%�$��0�����.�������������}�䢄�2]����z��r.�����~'�l�f8����ϫ����..�s�uaiW�O$��|kE_q���o>E+K�_z`X�}#GvST�R��&_d-<*SUnK�=ؖ��9vNx�)b�*o�ܢ�|P�ݩ��[��$�1>�q����/��@�*��]���-�o]	�nж����'AC��8�nh{I;Z��0���Ĉ��*��=���j�l�l�Ђ5�Dr���s�g$�vSU���������R�č�]��Dͨ}��L����?�bx�B��cy,P�Z�+��n0rd-J�沐�OC�u�lR�g)� �{
/F�?�!"��{��:���q_ǩ/AͶ7���ڕ}�bל@vI��˰�GA������a>�1}C����H��Ҥ��@,���'�8����Gb��D"�z"����m{������ˤ
����sI��CX�A~ﵝ9
�I�� �kT��?<�1�p�m�p$?ӂF2Wv5~^Z���-p�}滞+�4����<��oY�,\X��M�ާ��i RJ���Z��o�È�������*7��J��X�.�Qw�z��&�ޓd;<asu#I~\.L1�Tdk�V<=���w��)�9+{�����hz�4Ag��)����S$y�3ƻEE^<�,-���J�`�gd����*�7����n�)8ͨ�Ý4�)�|R��tV��CFت�sl�Gq�Z�W��w]��ss��Q��
�ı]�E�N��������u+ڲ�%�m�3J�0�2yT����"ϩq�oE�a�x@B��q��B��k}Lv����2�Ѹ�$Ĥ����d�j��}�פ�>F+��C�I+�+{��U��yR�W�	i�)t�f�� &����?��\�,ˤ�x��v=_tRy�IP)'�'�p�!I����E����'���4��0�M���.(��cAY:#���bW���K��&���QmGW59܊�_x��#+Oȶx���IC�_�2)�DǎM)�S�\�І��{j4LLj��p��]��5_�'q��ۗ���rt	�ޓ1kZ�:uN�K�w�ՄՖ�g�םuy7=��_��Qq
�=����z�:S9�͹%DW}��J�u>q����kvt�Â���)�uū�=�|�Rd��"��+Ӯ(�b��$��
�my��b!��>�X���DRK�Α��S�7��5l�c 7��Hl8�/L����
��N����K���ɗ�@�XW׆������ԃ�hd��B;HD[V�����y�Ʌ@�Έ��<Ə��\�o��� �Wn�4��|`{
�4�yW�����.��*0�&�K�n���Jz��}��'���8ɥ|=�?D8�#C܎����:a;P�Z"V\�0�[�\���Xs*�O�s�(��K�y����Dӊ&7��<dQXlX��bh��t� m�� �!�ל�}F�JΕ�b�35���
���uT�+ZߕТ-�&��"ae�X� � iЋ��O����Ʒ��?��/��g���7���/u�lI����}��	CG�<Zo��H��|��7h+��A���"
����M�c���N�>v$�q��6h�OȆ���F�q����U4��#y�+���3Z�E��?HdE��|���Te�/M�����ÄN��S��U�EP�Q"Z4�z�d �a��N�u��i<�$�ކ�^�ue�xN��I����k��+$x�I�o�z�~/��r��P� �"CG��T��bR�u8b>��<0�`�jR�������/��T����3ah�z���UC~��.J%�"t�@z��g���+o��[OU>�[��nގ���s�* �߃�����^y�xOE��X�9������X��l6��&��{����I�-��C�w��NAX�Ҡ5�d���SX\����tH��j�
&��*�]p�|�RϬ�J���#9[�/�m���`��j�g�Sb����Ѷ��n؋��Z��娸"+��F.����*��O'5񹅟lM5�;�.�>]��ǞRy��p;b����!(�V#�d��OD��Y�=�?����v)
 �O�ß���N�ۑ���a"����L$��@���}/���?)������r���疝�T���*�\զ����uo�G� ukp�e���ˀ�p�O���d��7� �7W��-T��S����Ѱ!��ȡF�דM}�e7�Z�(萄!~=��7��pr�)E�#�$�Z�a�	Vc�3AP��ミ�v�l*�W�_T����'X�����!2���^_��Z.9d���ttt�)�S�{j�ƫa�/�o��y�b*~Qc�!��y���t�����:	��hG�ł�<��f96�]�0>�;G��^��5�Q/�^1g�g��;�у�@Ō�������?79�8Ơ��^�>l\��{t�Vp ��P��uq�I%��q���l�Z�f"�ı�016�GM-1�\��&$��]���)�Y�Yۋ<�f���5e!m>%����V[(,:[4���+$�	z�|or�M;�_�]����WX�޳o��7�\�Aڊ
� mii�%L�/�ѓxHS33�$5ON�����W
|%ӧ'.��u�fk
��=HMꚞ��vE�=ZKBd�t
���v�D�P���%o��Z�:�hA�C�c�bh������!c����GG9�w��|������SJ�~U/���PAI��e�yI�S�������_lG��T!BlR="��!���Y	�M�b�w��C��̊�R������<��9ԇ.쇙��%U�x�?��;�5�=�VV�֏��%��\B }�/�&u��1H��{4t��olJ����Ň�D���C�39��q: WLEEE��� ��b~�`��UEF[���Pc��hes4_5�
^���d�'���aI
����T`�K����Qb<>�x���l���7��R����V"����q�/X�,H��C�B�Pm&�3F+�vo�]��;��m�R�9$-�^�UI$=��,�ٿG�<�g%��������1���Lff@x�8�����'�|����uĭ�T�����d�^���dRA��4���g-_`ä���RMmo� Ȓ�L	},%������xO@(�T�����5w�u���r5�����\A<]~�$���b��in���;5<�&=Wb͗����Z��q����˵�P�nHhD8���3�I�ײ���9�;9�)Mc�p��
 f�����FB���I�k����J&:����mn��᱓,v������9�?nz� ����$aZ	���U�ɤ�r���O�ؓI���plB�M��f�k����J��M �1���YV;;�:���չM0��&܃Z �I�Ā�;WK����(4��JGlb�Ǹu����5x�T��v-�7���-�ꄣ*+� �H\�d�n����2ɜ�������{/ǯc_=���~�>NI4���P2����K�<;���C���	QB��� �6�B�B��3כ���+�11�i?��!F-)�4	���
��s�9�j�/��OA\�W�����^�h���RR@�����vK�vj�^d8s3i�U^So۵�*������P�2o'C�4��	�S�+*ȅݍ��Z��7Nd��5�V��x�d�7CI'��Lfq�J��`G���9��JR>�nVwʋ��4)��4�V�>�	JV���ob<0^J܆`$�¯_1�Q���ܴ?��-*�$z�3����r��V!��V�b��;���#&\���ۘ�Vw��3�`�]טZY-�V�M�\�)M�-���
M���K�^�^]ˬ��9�x�����O)�Ra��wl�	��@�_I�x�}ذ�9���A�A� �^Tʤ~΃�)��6�a�S���H�F͌6z?ޮ��&*J2��Lq���sJ"V������VZz��4��]%����z��x�~ڨ�b�d��E`;�[:��̊=������'�挾�U�Q�W7��DE�gd�Z@��;��QPȲ��RＡ�����N�M�?�$�	&��������:6�L.N�xΏ��WsCNB�+�A��p��d轸�s������m��|�Cz�]�����W��g�zX��@�.�i�[���_������y�t�t���]�$1[R��X��<:�ڄ���L�߿�"B�v��&|B��Y+�����,j��<]	�ti�o��ޤB�#8��o8��硅� ��C��f*���!x
?]�̠�Lv��Zb�uZ@���{Tw��j#��=i2*���(�zudLMJ
⸑7A�K+������ݜ*���#�S-��r��x~{�� 4��x��}g��0��m����e�%�ˡIT�$�?Y_hi�y��"W��5�IȾI|��[��)�wF>P"4_���<#�~%p��6*�Q�L��y�Q����D�^�@F���Y3����V�L].�8Ė��kOn������i���4����|F�C1�/�U����e��`��ѝ�˜g�ҥ3QD��J�n���P���K3�Fa�Ս��J����K�~
���u�����(Y��Z�M���גX��f�d�������sx�2���:�퇭�AF�V}���TX�u�~����<'c����Æ�6�O������.�_N�^�Y���/�.ǅ�|��_s��4����xl���Y<'��x�?	��,8�#���[�qatݙw)�j�*OԚT06�"���z�{c3�+��m=�W6?���i���M<��8]���(��X@F��e`��{!��Qϓ+d��[�-���tg�Ⲯы&@�&Do��p��������4�X�*"t���q¢%L?���!�i�dmÈ�s��^ �����-q�N��Т��VfؙKK�]	H�A7�l���w<�.'E��A�W��ߐ6A
H���E��^�y��i�����-ZF2˯3?!HT�c�e�ۋ����[��?o�%D� �d��N��O�	�s|[��?*��N�^s3D�1��_�V���\]]��%I��ЁYm#t�{/p"�iM~}�&�=EY��<��c��xLȹ�eC�"��dCt7���*ĊeG�/;v�G��XS%	�=��I�&���@k���f� �T�d�9�u�j1�s�.+lG˶��.���4
=a�&+^G@�b(+.u����\*��r��#�QW������e�;k_ a�y~c%"#����Z��I����y�Qy]���]Yd��LY����W�i7�� �����-wiG.��Ͷ���@qL�Jf�	�c̝9�)R�vN{t4#�W�@mN�eKw\������j�ab�������������q��qTe���VE�
���X�u�Jaqd�C����[��
浝3~�>I��]?%@��nx̱���ɾN��Z����,�`V��wxP&�P���]F�yB�:ޕ��!�~�T����6��$��h�Z�/j�t�\�E��˶,�<��1M2��4Ϯ4��P���ܮ�M�[;l��|��t�~󟶴^�#��/q�{�e���.q���e7]�U��F�����c��<
��`,P�>��,�_p��2�\s�{���6�.��<D2 ���`���;6��~^��y�JR��&���]�J�o�޼��sq�3ع�#AX-�FJq>:�w��=j��;�#���#_.��UՖ���O�S�6fK��J�Qę�J��NES��@e�����,mk�&�{44�p�� ��ϕ��ԫU��Q�N��������?�itX��\�̙�o%L�8�Fk���8fyx��>"ZB44�����t�B�?��1\]�*#aoԼtۼ_�����}#\ 6-5Ǟ��x�r˖�a�N��VAU���'���XL{�Ql=0#`a���V� �	�.���`�?	l���2�����T�Г���!� AA+���)*c��&��܎od�+�eȉ�I	%��Ά�C1Ĝh߼�Q�t��D߼O<�L������VLa�����v��|�c����3��LTRv�Vf|�i?A|p���2����l������7P·uywVf��ΕmE	�Z����9a���/NN�C����G���#U<116`���E��(^W�����d�ؓ����m� M��L�C"5�˸,aU�F�P��F�����EY�4���a?�#v�B"��0�6��M�UP��w�M�{�{$�0��	1D�S!��˃��ۼ�B�uҾs�P݄X�Ԕ��'��ps5�%���-��uKU��ֺ�F��?5=]�� �`(�H�u��ޅX����Vub�~��pId��L�jiM�N��D�PR�;�X���*��E��]"�V &�<[ߧ#v�P �n�m�����6��ڞ���S��� aB_n���	�{�2����]��8��v���=��:�w���؇1��?��
�!*K[Jٔ�F��N淾j(w��
\ܵ�'�Ii��Ş�f�v���w��	>+%*Ǧ��M�+-��B��9��j�c�y�%`4,��}�GL��ﶪ���-�sGe+U8�QUF�ܧe$�{��
i�p%���'89�A��Q��)�Dqn)���=�J�7�{��u ��G��!� 6��M�W|.�tl���D���}�7@��Z����W����pZ�.6�*�0��J���Ǥ���>�^/�w��)`�{�,��1�MT��������:=Ԏ)���=h���p��l0q\��eŎ����g�jH�ܻ�h�W�M��J�����Jw\��!l��9#�?D$�]�.M ����ݓ��Ig&�=O�`�Q�����=Ws�>����R>n�>����jWN)���v��I�&Ia�h���x��}�+;�z��r���Z�����]JK�[K0(3���#�^���0ة�!p�ܸI��ʇ/�C ֜G"|� 8��qkv��Z�-�_X�8wcMGr��4xs����vZ1'���g]���L�v��s����ſx�D5�is__���FEx	l�����%[�o(�>�kL���,a��0 ^s�K�L���鹛&pR?-͢»|�x��� �x�����/���ց$x�?�zRVQ�[�S�)TY�#�^�M�Q���['��� �v��;�$y���:�@��a���0��pf�DG���z:j��/�����l\P�jIY�O2���B���������=kg���[?��q)�[�@��{�i=��mO4sJ'v� 	Z>V���#��,�B������vˍ��	o�{W/����aS.�$��\gk���?��Y�,ªM(*U|�	v4�G���x�eN��T����(#��SJkT���G����
�Sm3'���&��H�s[b���U�W�>��z���H&��\]��7��I���p��]]����6�s�gz���/(��R�Ҡ�J�L��%����E��t�'�s��'ӻ��j���Z��=��Tbw����T/��� +�Z2��z��2Pl�zA?|�zP���	��Ϧ��f����5��/�>9�nYZu�!~:��t�1D\�k�$K:;);/�;�ğ���iS��P�)Z5|
�[� ��O,}�m=�ʋ���S?�d�ɩ�����R��o�z��ś72)����<��*o~u����5`�z�s%+=S=>j`�5�"�`���jn�}_�T�4o���d��-��������f����	�EV�k�tj��iC"H���9�]S:Kh�R:~����PI���7��yE���[��W�L���h���{��|��Q�i�`�
\]S��x?�I` �	���g���O���kk7�l!�};�&Gs0� ���ݧ�v���\���S=��hVj0�"�����8w�8K$�˳!�*f=���.>�ng�g�2�#�#�8�cW֝��e�Q&�BZ{����K�xO��[/�^kRt;�Ly�_��"���uV�+.�g�ly*��58I�1.����w��C� b̟���(�P�n��~�zy{;]�j�����`+�"�vч��`ӥ�����!��tԫ�y��W@WC����z���b���yfw�����l�,�"4g��zV�"x--���E<�Q_^���2��)hO�[��i`x���ˏ\r������Ŀ/Pe�1Zc��[ê+�ۯF˧�*�S�N�������w�d�>.<p�O�T��m�9���a���Xp��걹�� �5Z���`JF������&�'8���/��e��Coi6g4T�aG��>�t����ue�BKK�G��e|���D����{�Xv��B�C
���Ԓ�K�����K�i�\\�N�����8f��Q��_3�M�F�N��ǹ�+J.%�����+~��.�IJјR"q�1�Q)��7�D�{���I7�^�mkRv!�\B9��q��?�V@���k�����>� ���Yqem�?,��}�y�B5r �`��ow�0��Ew���ٸ������F��;
����D��#�j�`I��B�	v���y��z�p��md�2|���F�*��x��=�:W���m]{ rd sg��\*�N�P�|�+�<y5��G�9w��Yv/��ͽ���ٵ.�����&�k�[.K��[����a������wR�����K�./G���a��
!4�~�j|]����IQ���]�?��5o�:�(�-~��"�uy�����\�L�v���#�eok+�]���h��~3��X�H�n69g�Hԫ�U��ӊk���/���� �7f2���� �Ru��Aߺ�H�A��I�)�2%M@��>GR�"`9�r�o�Ԍ8��W^*�:i�����G�zb�v�(�ǱT�K|�<F����s{��)DQFX��sX�7��Ae�#������J��?�v�����V�ݥ~�.�j����� ��ZZ"��������������Hao��-�#g�;�f���\�"V���q���m*�� ef�ޝ*�	�޲�ӕ��&Ð.+V�϶pap�W���'�Z����i[�F�=�n+[�T2�t���{��@daaA��6[�%pT^�k��a�:����B����͘���e��ӓ�F���c�x�Bu����=���66(IIIH�/��O�iu;�v��3:����egl@e��7ajGs��&g�f����Ɏ2DI��)�U�+�g�a�7��L��'B���>�(I1%��dK���?"Ȁ�.�!��80�I�d]��w=�b|}�]�^Xs�g�o�TN�D<==}�!|R33��dD(����� .	�Ŷ��S�&E:��|v��P��z���l@�UuR����sI�D�vo<V�C$V�)Ĝ+�h2iiݮ����30�����|���|�l��6��ym��.)Dǹ.�3v�!��h��Q=��͇=�H��;�î�������lX���O�[ii���bϜ�A�����,AV,��RH�4ɠ���T�#.�5��l�t4��g;��%͹�{|<ZK����*��f߭�%e��۟F��o�������p��|�n���PI��e�z��F�>W4��~\���&kvÆ� � tI���D�w�����k�4��;s��"k���qk[ی��B�.���4.v��*~���4�R
7_)�h����u�-gb��
�.?I�^�}�b{�t�GSF��H
�X�齴���(�Z�C��3���pZ�ĭ�Ϳ*���� 	�	�$���E�Q�P�Gt`�\�%ГC�F�u�WE�5�MCf� W	��\�e��Y�F/UB,�tF��TG���(X98��������㊦5g�e�0¥��&��|e���z����T!֢��� �VW����s��t�џn9˰�GSǨP�UX:״�8���	 VQ�-�.1�,�g�8�aT��8>�^[f���|hS��3�=�ݕlл��锎�F���S�̟U�2���$M�A���d��;�Bu�B����%�|
���&�él�/�ٺBpŹD��@�ws��D���3S"�P�&v7�[,�?�<SKK���IM�&n8+X����T|�Q�p��V�����O���T��Ps�x����2qC�ޜ� �pH/?4q���
yy�>�$#�1�4�?M0�A�G��������D#�OFŀ<�^ݰm$gb; �/4(�JH���	�ԧ�+�&�Mx2�i�(�I��Hf�Is�=׻��/!���R	_i�?ije}��|wi M��HVv���iٸE濡����-((��R������V���%%didX�e��	W5������͈�vѭ��e����d�ʐ����&L���" 	^��dĉE���.�P�c���z��u�_ڻ�$�*�4�ת�C�\V���@0�x*����l!�4<�8��m="\��Y�a�#U]�� _�,�W'oyɰ�9u�OP&�X�r�4N��[�Z�+��L�k�RA�1�o^E�ߔS�b�:�*��{�g#9#w�*�^� Q�RT��L��:P]C���+�mN���Ϟu��KJ�)��
X��	��y?H���7m\"�b��?v���Y؋��PT��Vz���%��' ^}��bk��|U��(��$�f���$4�wdN�ΘW�SU�o���ys�{zM��Dl>D	0m�U�L.�g��c��ܻ�'��M4���ρt���(<�jL�;���0S[�enӑPzm���NW��w���g"�kM�K�9����Ză\/"ꡨ(���x߷���Ծ�Z[E��e�����{]Ws^���p��TE3B��	T��{�۲�5���t�A-4r%��5�Q�{����_��5��ݼ5�6'����nʕ)+O���b�ALփ��-.��\�� �~�����a/���A`���q4�,��@º����w"fSIs�G�99}�_��[7I<Vc�h��7���DZ�E�;��*r�q��9i$4v���a�f3c ��?@B���yG��^�=��e������_���f��D��Z��sE��dBL��z�o��J��;���ݏ��F����zT��G��k}�f����W�;��玻K��r!�f���Ye*ש{�M�N	D#VYÙ��P�hi!)�b5�w��N�K槢�"��NZs���Z~�fδ&�.��H���*Or�b'��=�q��6JE,�)�/�x��w�MDI9x{뱶���ѨIw�wU�%�q��|����/���!c��-���}m��S��<_ٳ_�6�D�G\C�K�S����<�ϭ���z�������7����G��=w�p�������	�Lu�32_iI����'{{�sx�Y�[���"��)���<���jl�.��=�YR�5�V؄�eSx�P#C���"�iO�=���*HjԴ6���͡QI:�z���j��בA�5�^��-�Ѩj8�zgfX�3{~6 ���:q�N���%=~�|M�/ڪg���=t�E/�&$���G7�4����T^$$�:(�X $46^�;��7v�w>/sϷ/�h���
�B����ݝ`o<�w��۳�Z�8�90Ŝ�MT�AಚU�����z�q9�uݲ�{}tŲWr�K�-�R��{wk3__�$\�fknn�V�
\H�� ^��ɹ܄��%)[�ğֳ�uK3�@j��Ï6O�ô.)�׎�\�X�Hp"W3�o:s��
y���=���P8��}�;: ��k�X�����BB��>5D���V�B��#� *�&�[$�&��O�	��-�J���E�|}��]#]$�y�$1�t��I�*���%��c,��h��-�����5�D(�]D�2��An���O�/���_�gg��#��c5�!���p�eB��m�QI�����Raj؇Aa� Ŷǋ�ۋ��L0���M{�����r8�L�����v�Su�Rx���c��HFoZ��j��2�7j��-��UO$�_v<�.VLj��j�P�)�d�t����$KL�k��7�U;Sw/�$mK'7���(+�o49���%m��f�$h!~�'����֥�H�@��-���Hm�f'��EuOH�,���ӳ�l�z�̮=�A��W�x!����vg����f�7t�'y�?��B��a�a@q�� ����VK�-m0V|�[x)����u-���Dd��w�/�dfv	9�|_&� 0ϕw-�pJ�p��M����0��N�Q���K��k}�${g��at��Z�$��;��c_v$Ђ�t�ܓ��$J@�/��+��QW����vF�s���(��Vr�� �	a�yS،�-,�C���\�Q���݁hs��K�u/��Jk�e����7sB�2�B�~a��{�̮�~d�o]����$���_��Ё��zY��gy!�,�%/���dw�����{o�����Z.rOE�<o�[Wo�#�ycU�-��R�Sr&�/����q� �V�"��8���&|v�S���!x���NV^��z`��w}�G�Іث	��}�IY,i({�~�cK
����P!Iy���7���+7@�FfQn�d�@������/�BZ�3R{���c�7�e�Ys��߯�c@���J���ђ�$�ۣL�ɽ]�|�8��Nh{!�o�r�MC��G�K��)E���Nn�@"v�6��{8�3%���0�}�E���Z �:��v��K��R2�1YvWp;���_n��7�b+�n��z�Z.N�EADH�{�����q�.��M�j�����k���=�U*�]�����̡[�ԟyM5��i)�%��t�n)��+)�s��R����6���!޷_ֵ��lg︣~����q���^ή��75_S���G/�V�`�+��.gv�%���}{�[9x% p컰�Wkfo*�YoH����T�@%V�*qNO��+��@5���*��}�3h$Wt���;΂�� @*�}48�CM�H���C�K0U��=E��ZZS�9�=	�\����z����O�W'V�l�.q�n�S��������nE�J�K�{lCO���y{�>�/���6Zf�t ~-���'��X�;��;�,�[qqp_�D��U�0s��YAV�j�����+�W%ϕ�M��w-w9�<Q4R��9�1!��l��7 ����KXg�9��l��S���>ׄ���ŐҤ(�|"1��<���b��^W�/�h����0xȀY��ۛ����9t��	R#�Zΰw��㒊���(��7�M�iS�AK1��3 ^�ʋ\��y�Ӵ���R�g����:>�1Ek��,	�vADbmT��.S�>��c��X�Wu���S����%I�_�#�\,Q��X�����Qn?'��,l���u2m�LS�Y��R~�:	�|�.^U����@.q����jK|Ι-�h������M�A���,Mz��-�X(4����U d���ͤR���]��\�U#�Lz�����'��	^�&�e3àN��k�\�88���A���u�P��z��₄�����b�ǽ�Y.��7���@;�c�M�5�y��֡��ϙ�
��W�LW��κ̼Vn��R)�PB/r��K$�`p��(�9�q�AQ����.P۠�1k�u��.hf�F�4���9��U٘�6�|5� ��W�$JnN�7�,j}�b��sG7�^	�\&�Y�`X=�������z&�(�Y ��@w��K=W�"8
_���_�"�1�q�P�ݢ'�c+����Ȓ�-d���	�B��f񃃮[A���6*��;j��2�%�����.z-��w�ys���-���a����cacۂ]�7�{�jS<�ǃ��6gpW��[=M�?=ܘ�١��}d��t*J��ʍ����mo���p��J|���f˂|����c�`.�m���9��8�$ʍ�'��m0��*ML��V�9�O������C�m�����X�ؚ�M�m!~�+�_�R���B ����^x��	���������X�a`�%7��O_�;U&�{h�RLa�<�,��iMu�T	D�Hi���B�*��Y�2p$��A&��=8��R��g}>�eY�\��[����K�Sa���.���І	���c@a�I��RK��FN�`G�h���}�?��?V�ƒߡs����9�e�8\������� �^��ECj�ΛلH+���\����֮I��&��-�{A��+����X������9�;�o��)�Bz�no��A��
>�f�R��ð�ȮHF~�X�v4�6�!����p7i�񾱕�R|u�>1Df�ҟ���KT�(�T�>x:�ෟ�#jL�+�z�#��2�Ǜ��2�jT^P�v�$��52uȭ�͋\�D�GP�z[h��qev��l���d,�h��u]jV�Oݘa%"(����۱�G%��jЩ3ҁ�Hπh}u�P �����|��}�9��N��u+���
�t�,�ގ�����OjF}3;�po݀��+�7	5ؚ��|���s����
:T�*>�խM�Z�.%�"Au܂��f7����
�(ϾI+2�F���R.>h Ƴ�'$��y���l0����G���[V��1H�!7_���� @x�`�`44�����ɋ':v�r����;Z�!r�`�u��s�f���Q��8�Y�d��,�r�m�Df�D$��-?Ő$��e�jb�*�������HGn���Ş薢�k��T
b3�P�g�5wȸ�A�����c0Mw�g��#�����
 �3��Zڢ�_���,�=ab@"�f�G��?�ڸ:Q�v������ORN��:��O���/ֿ�G�q.��j!:�أ�#T6�X���'l��H��+�C�(��5;��t̤�L�=�w�-\�.��� +�����M����g��ԇ7�s#���B�j5X�h ��4b���I�c��l�H �Kzی��Cɡ�>
(�t �å�YY�/>q<������Ah����۶���BH�h���'�,�DTI��MZ���+R/�,'�G�SS�`4�Yܫ�+�� �1�����?��3��ץ�����9O�)"���b��\�s�$�:��:�B؍M_�7�����O�k`3a����zO�ֳa��S�z6���,u504ƾ�۸���c^�c�� =�����*7�fb�4�`��y�>�DL�������}K�-Of�jNA�D����ù:C?I�X��/-�w���ޤ��n)5d���˷a~��}�I��?/{�h� Re��°��:�#%�߳0A�o�_��c7r�ܷ�0��W�
�o�f�R��W���yX/���H�{T�I}���O!�@���� ��~��5�gq�������i%��z�ǉ�.�?۷�1;
�3�&�R���TN΀���ξ��0 �ᰄn�c�@²��[@K1 ���߆�t�/��,F�X��]� ���r����b2���!1�}��xfV�v6k�D�~\�J�<���C2�S�r�D�d6�+�u�uƘ�h�t�$�(�	���{-��I���̝�Ed�BC�Fw#���)`F���U���E20·O��(o�|R|#V����+}s2�}�1�Yr�q)h������$Z�Nz���Ƹ�|@�U���ɣ/�Y��	���g=�a5wd5��O�^yF37�6�*usr��?��z� ��C�[�OƖW/�DAj���1�4�Y!��ט?!_�`�Y7Mj���m� ,��75��������wf�<ޯ��}�-고B����r�P��d�Rw�C]d�Ć8糛L,Q~4}Q��ko����{���F:4SkA�UXa.�3wgْǊ��U�yA�Wͯr�řFoX�Z:
,���8��"��U�&& l߿ T�-��V0�Ǆ�Z��]�Q�H23�UHJn����������g0��?�F�D�GBD�F/�;!Q��X��hQ5��Y���DD]m����,���g�;3��1�b�\�U>���>J[�h_�N�}~�1N�H7�܁0�0_�@Ρd��P�ٔ8C?������k�2L�v�lۂl�B���<���u�Ϥ%�n�4n�������b�]Ip��7�"���LJ�C���4hu�EB(���By��{TG2����9�R�n���������'Ŀ�sGt6s����nt��qT�=-x����Tz�"���Vɫr.C��*��c"=uA:MA��`V������BA�-�
�T�ӓ�k(wM��R�K�:p,̢^罧�àT8���[H���TF����<m?�w_��k�b��n�%�Q��Z�0�P��l�i�a����2�N�֎w��.��B�#
��@k8!j�Q�~>[~�d`r�^����A��`�k��SCO������3���7݄�J�|�m���MXfC��)�ꨋ�Bf�i�6�?d	��l��'⹁�&w �t��5�?��:M�k�tn�w,3�ds`�?!�}�C��nr����|Ww���"��X���jgz��o�c���=�'������j\c�!��3��>�����N��F��tn��.�bO��5ު)�9�n��Z��ǲ̪T�.���*�&�	fi�����.-�8?\o�ރ�#T*)<��W~1�<�ٙ�xFDo��~
�
7R�-{�����%u��}u6�$�2��#�-�sv�Su��ֆ\�\��\if��A_音���zXp*x3�4�A�I���>���u�&H�4��|N������ܯS�R�� t�c��,H_E���%��擰�?b.�J�������G��:w��]�w��6:3�9��t�R�/t̝�W'#,D۫�]��V䕬�v����<ڧ�R�PC�zŀ�p�"��ow^�Z�7�&u�R��o�����n�6s5BEo~�MW�rdA�+�4*��G����]_9��։�����S	�_J|㪷����B�0^�F�
�D����;,;[�VyU�xeL��e��]� �͑�H�\
}�aϣ~J9��̄����{��L�O��Q�����x*
b+��i�<�&�3�<����%E��i���W߼�(�]�U�����}�{�$�aQ<�y�x���)J	����g�X{|�ڪ�{M�S+�^1s�ڨؼ#���o���Q�3&��G䛱�L���tR��رg���_r�Sov?L�Q���|��U�Տ4�CL��U�mx��!�˨��T�ų��A�k��@�/wO��T(lt����;�����E-//�L�=S��銨e�\����<��Ǘ2�y�X��'��u�IĪ#�b$�T w�'=��uV��I:Zx�a�u�u}W+i���/�O���@:	@�����(x\�H��[l��61��ծt��.�I��>sX�;>�s�(���^r�HU�8b�s�D����.���|'m˗#J��yX@��>�:��$���Oij�O_�r�S��5^|pu4��Mm�fS2����R���T�wȚ}���>a���Ѹ:t�l�p��2O���qR,k�k��P㚮w�%�ٝn�G�	�Yk�5��>b)R�F��\�%O��v�N�Ot�p&lt^Z�����~3r���6m�4J�U� �g	/)��E=���o����2j��-J�x����ۺ)��ц\�`X�j�nUjdr�U��;��/���!��3�yo�y�}վ���>��
,�l����d�bV�(�F��ԧ�#�Zǧ���=�vMvY&�/:���8����X�[ N��:����]�������<���b�{n�s.���1�w��������R���$�ohJY�v0����>.)��lp�M�xw��?���, (H�W�h(��� 6�Nl+����h���8^��{�p�������'	Y��2��5K��;�	�C �=�?�Y�d�fhu8�n�U�"���ba���Σ���K���q����;]|�&��eG��؃A �9��t3��9GwAwEvVϾno���Ci ��w�_�^w�yƁ��;˧����	��XH(�'1N�f�\���k�-60Z��m�:QtCf����:�)��_-0N���-R��8��P�x�u�"��s	�"�wg��+�z0u>`��~�����r���G�X����)6�?�[���L-��w���&9�l��ܟ��a�����+d�$����u	6�¿���c+��pR0<ɩM����[�˕y�?͂4��H�c�K����L��\R����ۻ5��4Yka!]�R�l!��1��~�����tQo�)D��#�,�h�0P�Vo{��UǑ[>v+���:�R��*���XʟR%���ν5%x���p�
Z-L��~�u�2W���{�m�֑�go>��;�[�2G83�t&���P�������Qҧ!*>c�r�]���lb <�L�ۋ�p����^�4Q�J�5��_�U�u�L�֔C)e�zK?��]�>]����ߠ��Q|敱���y:��:��Σ_���\� D��)��XU�~�r��I���_jRX^p4(7t��P�5��������X��*tg(X((L��� C7�t��U�=N��떬>���e��5�b�jo�6��je��J~���v���C�4�yJ�󤭒GJ�,/}-����$�,���-����Tͧ�И|�*.�S��j�*�&LYn_����+���� ѯ���וB�M���`��P���e�}�zm�J}�[;�c��܋�($�1~[O��(��ڛg:TXu0�	�t��\W�0�.�tvq!�|K�zG{..��r~�����M%���|��ܦR'1C��70!p�.A���,�V����}��J��~���ޑ[q���' �8�S���S�:^X%��f����ݛ����`�p:�Ic=O��gȲ+3�m��r@�ytJa���%o�E�����Z�څ�~d�h�,������"�DOyyQf 
��������P5ZF�����߾}�J
���LP�B@ͻ�3��/C^Ն���H	�`�[5���l9c�K��G����Y� �o7k!�6���y����jЁ^�)��P͐�Sf�X�C��a����<k��|I-��'��KK�ݽ�8�<ai��u�71A�)���oi�����3͆�ZRtK��K4-:%o_ }Z9�q����vԥ� [�����'m��s"\�B��sp�^��!1Ch�3<Y�`�j]������T0Kna\陠1�#��ܽrK�C��:��9��'FC' ���N����	L1>�Q*���t���$]>��ޞ{v��/�b��c�3��Z�"�5樼��t���&��z�3�#so�\� ���'�8��3�W50fh��^n/LW���\"P{>C�Թљ�CW ���چ���Ӻ=|^����ķ��la���{忘,!yX �
��(�i��GF{vU��� ETzϭت-���f'AD�N$�J�t��+A?Q9}�]�M&�k�����t9�4<�a�O&`����z����Ɇ����Mi�����թ��_mQռR����&�_��¯����e
T�����JdN���_>�Nِ26I�E���͉��������П��i���+�|Ȝ��.q��(�[�oZ�U���m?���O
�e�_B����p�]#���N�n4�r��#IA��-�Z�{gm"is ��+1̴[
��ESi���h6���=���m�޴^�U�"��j�!����p{�Y����S���^Tjo�&W�� �{6Re0m�:�ۍ<۽1����Մ��rB*s8)���b����)���� ::�[�BRe�2��ن��G�%�OI%�a�T���MF�>GCšf['�T��ݛ ��fA��o��x�� \]ŷ?緓��O>�Į^����S%�lWIS�<8�U1��y���/M^� �t�������kA2�ZL�Թk�k͠(6��QV�o/T>�y�Aa=.sI�sx��oK�P��#@��{N��,c�QX���~b"���_qϦ���*%d돲�̣�	��+5���<��֏ף�5��s�N2�ƪz//jɶ��[��½o
˄Uo��V]��DC��z��}�-\��=�4�h�m�I�E)i�Ypq%>~A�Hv����x�� W4�<��}����Z��p��g��n;Kۓ��Ab�TzD�!�w�/�1HG"��ln����P-(�.(����Ӹ��)eJ���;u�(��vV�>�_�Z�0���[�O�G���Vt�|b�R]� S2�c�#�኿�є���~b����Ϯ��/�a��h��T��N�<�Z�E�R'�Y:D/8�R��K3Lj�"��<��/2'�����tyN��0§UbU��#J����11�RbD%����eM��~-�m� �����Ԣ\���zA	��Q�~�f��귫Ӭ����A5v�e�#%p��k��RU[	����sJeE9�Σҁ�hZ�#��x�;L*�����Q�յL]}�s	��b��q'Ά�S��F_,h3�qid�n4��!{���/b ���QA��c�Ϟ#fEJ���N7R�~쾤��V�����z|38���a����u����)�A�m���ש�JW+5�lw��Y]#�~�Z�<dF��k������TA��M�Ѯ̯n�E�w8�43�}���.�� l�=_B���e�8�B��}����*8�$V*R\`	�<��z�t:��<l~�tV��#����+sȟ�-F�!��!�ŜPO�N�7�Km�����<G�lд��.p����)W��ǌdXm���[$�t�{ˌ�)�KT�ֈ:�h�*I���f�i��T<ňd��핡*�������g����87dV��°����J;�k���w_�\Y �u���Q��ed(zg�PY��oiZ��d����4�v��""���h"�ީ��1�@��_��Į㆜�w�H�ޟ��2;OL�}�o���ht���4���@l,߸h�no��Q'�v	�ȼ�-�!�WվO�E!��<�#��#��Q::��>.~�@Fgrtyo' �])�����v"N? �����MT�V���,�L9T��=��d4�?G��6P��x]>\dpA��M�&����bه)V��܉M�����u�;
=->�ubK�V����%[4�]����Y�G�}�m|g��N�5~`��f�ѿ)�=�������֛m��71�:��������-�vOͥ�{�?���FI 	�a���Q�j�[:�r�az�wҽb�W��ݢX|�)V�v�}o�1c����'������ �@n��϶9�z�[E�9W�T�UQ]�S���!��p3YT܉Zf,�&r�V�-3�������v�X?�l{A�+U�p:?'z�өCE�Ot�2��F���E-�G���v�"n��)L�������� {�w�e_Y-��W�"�x���`Yy�d�.y����}�޴m����f�o��N�����+�>����RD+���f{(��l�-}�j�V�j��j�|�@�%�C��d�x����Bk �<s��0
H�gJ������y�q�8e>��6<��$ ��TA0I�B3T�'@`.0��-[��0h:��q �{Q�g&w�� |B|��[k/�[�Ns<�{��ޓ>�yZ��c!H�ƫ�^CC�����{���Ñ@���~���cG6�f�ʘ���v��Z���!��#J%\�p��������Ǿ+v�m�|2Ǖէ�8�2:�<�99���{]�J��ͶD2�%�j�RZ�Q������/"�c3T�Y(ZW�LCѠ��'�ʦ�s�v��2�~a�o��|�[�ywK�NK5H=��X[��Fo�ڿ�`� �i�#D%T@����ŏ�K# �j�_�G�n<
K�)��A&@ �Ā(!�%�GG�oض:��N�~j��篐���{����i��s0B3H��ī���z�/mwq���Be�
I?��L��/L���fۈ�O��,�\�-�J,V6l+�*�3�0����܉*���L��h��y�pߧ9F��A<󡻈["� �]�6�@���=G(�OMN ��yc�=	-�8�\�.��R�V���7��Ȃ4G]ir�Jc_ξ_�SR�*pm|1�>�5��T�m��kW�Z:�z����3R`�#vZ㢔�ɐ,e�X���.��O�ͼ�0q�������KB;�x���_���˷�ש�㋱^���k������ ��O�HN�C������>����ӟ�/�N=>�zC�qM��ڜp	I��v����V}��[�k��AJ���e�|��25d/�Q�+��	rC��'[����}�[�*�O�a|�>\h�z��[Wl��o>�
��ncSFj7I������_y��Z?j9\f��|�3��E�A�L��~��#l�tF��W
V��o�I(5��Pm��P�/+���-�+�k։o����/N'm��1��?6�#{��@,�vF���6��R!-��IJ.L���B%��� (X�ԌL��k�f�hgJ�Ҳ���QL��<��~&R��}����	oZ^����SW���B���R#z /��"$��u��R
�S���JO�t�v<�P"�-a���j\�,{8�=Εd�B΅.�O	c���,��	u�����o������z�(͗�#��)kb�W����e��.���~ Aӣ���r\��m�j�v ۥV��Z�+3�����q�y���e7\��Z�2�%=�
�j���^�&��Y�����"�C5&�Ǹ����4T�X�Ð,U��0�5�W��v��J� �wjj�����+{��Q�;���`����z85>i ���L���Z�Nqe��Hk���Tqx��`C|�����=�D�3	�ylE@�-�S6�����C����|�ܞ�R*�:���~Va�?onC	dn@�����Dk�3�s��R?��4��gU��e���]:�ѧ-m�
qDJ�,Ќ��s�/��0o�?j|"�Һ'D#�d'i��0(��/lyݦ����7�ۦ��$�1'2O׃�&��~���&U�nOB���'ˉtg�����NBT�u�G�Zҗl����C�Q�U�Q�� �{$��O���]�Oko��؝5���>_�� _��-�04�Z�tJt���W��nB�~�e�]O��G(	����$G�U eR�y�xOѻ�y��.�4E}��I�<��Ҝ���:<���{!a�$
�}�����)^�8X���aa(�z��T�cPzQפ�bw���>���^�Y�͍,�����<��;�|������>$E�m�b.�-JTJl��0Ԕ5md~�ܣ�,3�D��:�w �ȗ�_�6�+���8���q�*X������"8&-�2��^jW`�YR��T�8]����F�Z@����G&�R*u�?�or8�J
�blr;Mʴ���A���/���lPi���D���.�0��'����78q���/Z��0�z�y��mT{:��H�{��C7֐��1�����Ṫ�� �<��W��Rρ���gX���->s��I�s�A)��/SX���8ӫ�o�(D[�P�����MW�j�
��+{~ciu싈�u��������w��^w b�V5`Xѱ{=}�Yi�~*��S�ļp�ދו���C8��]:Aő�[�F�ߧ{�F���[kۡ�TWR)Kj1���}έ�?3�G�����ⷻ��mY��̡S���9	�VO���BǇ���RP�N�.��ԙ�e��6�8���g�ۇ�﯐NSD���zw��@/Z������/�RՋbIR��a��1a�v+K���'�q��;�"%��
K�L��[ȋm�8���+�R �"wZk��'��kq��{��m�a�f��9��涂��ߨ���SԦ_�.�P�*��2�a
����zw���f��8�b���q$8���$^��3s6aC���-�F�v�T����O�W�"��.'�s>�v��Q�ٳ��IyF������,���sqӢ��]A���i>$��ű��eΐ՞�ձ��m)�*��4�	> ��N���<�~��\BO��MF�Y6��ƨB��_"jU��ju�c�m��u~���L1����ǡ��$�U��ᦦJ~v�DlgCE��%��V(�H{��n��='��>�׾A�AQ�Y����7�٣�wi��xX�����1y�{�'����r�����-��mEom*���?&&sK�ڼ:�$�v�l�~��iF$n��sGj]O�%�����S�~V�z1��h������?�j�nRm|�ϓ���KϺً�,�Gx�+;Z	 �\�q��'����[fק��,�6�6eu��k'�v��������=�9wcY�K,2HL �+u6�e���{�~Q<����J�؏�p��������N���#���;�����Г?a��z�wB��K����:�2�`�D�l�A}׶�{�^�㬫���S�~b���ч2��$�/Ѧ�?L�'؅�N����B�P1��/�s�s���ƚ��� � �/�(���+�l9��L4���Ԓ��ґA>�
v��<7e���Դ��`WI�`�$���O�2E��ߒ�/�W����'/��8��l�6L-?�U�D#7��!6�>�T�>�,ԜM�b�J��'���8�� ��5".~&��я���E�;�ÿ:R���=p��>��_n3<�H��z?"���p��`�������|�U|Ѳ"1���fF�'jk�~ <���!]�y��qLW�*��n�����PV��!��=ɤ�K���K�y�S�g(��	J��L�l��GŅ��e�q�;C�wWV	�����:�4S���l����`��+V3_�U
%$f�^H8}��,�e~S0�Y�pdZ�����wpfW�%M�X�F��q �<�:�,�a��i>��	�]i�`58��fJ��:��_p��ȸ��.���+F�)�~kj��w�;�ʬ��I�L��-��hf�]�(�f�xBƨ֮@�9bG���;ag��PH;�G��=�'.)$��Y��|���n���0/g}��D���:�4�.ȶ2/� Y���gc;ߜ�B�����疐�PX��j��En��@��R�: ������:v|�����\�N�������m���4�����a����Z?�ػ�SZǐ}����_|0�U�Q��w�䖀J���}�}	;K���mo��O@�H���=w�Y��P��O�~��E-<�Oz�W�N����cg�L|?����J�U�u������gb)~�>�k=���5Ii9]��DW�sI��ݴ��[�$�?�m�X-��_+q����m=��+h����������� >fT�}2��({�[gs�[���8��m|���l�&<����F�����'��S�����<���n9�O�����z\�$hn+�j��g�Z�F�
,<��HA�$Q��DVrߍj;��`L�x��4ݽV��;����[j񚉌$7؝������TYE,��4���z���R
|�@�i<�3w�7����P�S��9|�l��e57٢6�c�Q[5�S�<Ϲ�2=���<i2� �\�>-��h;���,�H�i�t�b�X��q�6�ANf~�$X���,��uJ��o���h��=��3��+�}�t���v</���5W?|����J9�u�k@��nb�볘���u�uh�d�xV&~Mx�V;�N�6�P6ӶDCc��;`�� r�ſ��|ڴ��E��K�ULym^�K��yW�B�m����.�k5��&F#�i�|���.��n��>��;S�TVa�#�KI�%l���b��ي�Atз'P�
@�u���⯐ƕ�z58[����z���UB�%�)��仺m�Q�ݵ���
*�&���C��$	%�`W���5H~4�cɜ�P���e��6��ۤ//�t�!*������e�	E�ox^p��m<OQ�7�)�;��%l�6Zۋ��o����w�a��ǈQ�=#К�����0�x� H����� CLG�¬K̅l�y"Y���٩�yT�,6雉�؛��!�r:NO�8!�y��fF��#�5���������<B]��$�xC�P=}�
#��LMg)Z�s�y�MqA���l54T��n�Զ1$�o��П��xMI0=������&�|�1�a����D)�X��o]ۧ}����$;/��r� ���I�"6���ȸ����Fx�2s]T�de��A��[k���������ȣ�w�5��)�M��V�A�X�}���}
>��hv3H��o ;�<	d��;����v��Kߪm��X�Nf�שWrYs]o*22�:(Q!2��$v�ןmH�\vt����z7�j�՘eY匞��p��%66� 2+&;@K��ƼY���(~��QM��Ae�7J�PC{vLl��ͺ�I)���12x�9 /��M��SB��Suy*����fC3���5�ic�?u	g���V��9�B�DM����<~�$�X��qU$�᪨���:㢽�$;��G�S`Z�%Vs���ky�&�k�̀�o'�J�9���E{��_�S�π�TD�o:�$����Bi�_��4[P�T���{1�T��J*=R����^�B��r�5�H�Id�Eې�o[�a[-[ʣ�B�w5��7��q�;=���;�r��[7M3���!c�6�j_�� 2���l*[�s�;Aͮ<�UX�ʨ㛥&�+���{6��C[N'?
?��2.|Z�`n�m��L���V�@��86���O�mQ�ę��!���W�=���V�ޣb!-�G�-�W�X�)�(ܗC�l	x�(�������}�ݯH|�jK�i��K*����{��a�.��+�W� Kk�����%b��}����(e��\W�TY�����=�b2�v��~)�{m�;m;|��m«,���\|����8��jy�IǢ��lͳ{E��r�7���uw}��1 Hζ6��;X�~Ѳ|7XDJ�*��R���{�[����X�y1!~6���_X7/�t.5Qު�y��(�5����"�)���Ao�\�u%��X�d�DI,���/Z|�'ַ?U}�t�I��<ӱ��qG\_4߳(�?z,�.X�G]�G�����Id�B(��r} �c�6�r/hl���(��	ɣ�3�)`�<�Ӡ�������z��>��S�<$kya����X���\ϑ�1���^��Q�]>���°
�|I��6F�K��d6��F�%�>mX"��(M&�[�A���Y�^a ��wy����܂)�s½Q�iM�� !]Mғci�O����MTVYx�{ζ��u��MI��ؒ��Ԕ�ٮˢG�F3��H��)֊#0�O�s��}����X]S'�2��f��r�$v�c4:OJ��/C�s�i�I�/T�����U��t�I����1"I3�EHd��T��C�6�x��"��OSt&��ReU'�����m<�ȼJ܋X�Қ�K�q��|�o"��.t�D�B�v�*r��P��X�G���w����o:�o �V���l�6�i��^i�O���@Ԑ�?ΞoU��|�j��˥=8�~�䇹�!��⊧�5�yL�]z2���u��X`)|�4Ų�
�!��cQO�j+2b���U<�X7���f�0,8�~1t��/�1�<�/��h�v�iM��촬�ό�10�r�5&c�xS��ޮ�U��E��Z2�b���1efoO|-/ʐ��P��ȷJT��/xO�ط�����꒑l�B��}�/��d��ҏ�Of�rE3J1�����[�Ǩެ"��t�c�>Y���~j�j���F��X�{`Ù%�Ĵz%
追�,��T����@0:�C�+��.��72�����яaC�)�#�L�ʳ��J�r	hkW��O��މ���f욇�%�T�&g2��QE�9�)ڽ��}��P�a*���~�M��J�9��7��
�t���)$0�i��6{D�@�����i�&A~!�K�I�Q��1����M����cA�L�6�6g<�b�J�Ĵ��<�*��B�hj��ű٦H��{M���Q����l��C�%^n�L
��HI	�Fc4=�L2^�G2���Z�b,@�����=]b]"QY��}�_Z�ZC6���$\�q�,�
C��ҽ(��Cp*ŞҸ1��r����<����Euӈ'�����VYhZ��}*�[�
�~��?[�˓I�?�fK*>�I�,q�iK�!Ξ�l#R�n#H�U]|A�c�1��K��!��M�O��X�d~���r��2/�qoП^F��&�;}����	���<����I�&KތT���ድ&))r��Ihm�i������)�� c��k+\�{\�gٟo�S�I-mE�J]�9�\�ӭt�T��CX��A-�㏞Q�-�������[
�IitE��p_GeE��+t�Vj&��P��|#�;��6a��}���-���(�E��n���}ޮ��>�P�H?s��܃���m��3W�����$c�F��`�َ�b���]X��k>�u>�h&]lS�>���'b��b���Zx�d>�%��1w/0��TZrw�o:�_vt��4J=���ͭK�4��>Y6� ��[���/!6g��� #*���	�`x�2!v��b8�t�K�����;�����k�O$����(���NUdh�('�
�\�������(�:q��� �g�|e�W, (EC�)�Ak����v1��͖]H.�1�q+!`{�_�����-PV�at�R���c�q>��)��xv/��l���]4�/��ZN�E��h�%1�m?]���-j�s.&��E�:�--���]�=�,�V_��8�����3�����^b�T�`�4e���}�g)��}�7ٸԊ���9�ekQ�n
;o~W	:����~��=Q��!���nE`�������}��TI��N);З�Ђ��nN�v��������S��:�:�X3�z{ͅk{G��3��X��$;���)�3+��Ԟ�d���{Io��+�M|[��U�*y��Ѝ- ��!!I(��&���j�C5QMf4�|-Y��]�j���&��8`Sf���-`��#��{kmI�DͶ6��D@����e�c������i��s���S��wN5�::�kV�C��B��G�f��}0�VL4��p���]H��w�հ��a�&����}_/��ꏯ�*s��m���H���&�<�<(!=�D{T����汆ݍ���y����$��z��Cz�:?b�Wά�2Mx��c����|յ�۲��үN�mY�Ԟ�Ze�p������3�_�]�֘�6�ָ�Bw�
?F��;ᔑ�7�,���kb�ě�9H���פ�@�5V��KJ�reIt�v}]�CoED�yV����$H+��FDD�Vv	�9�j���X��h�99�V��$�y�{�Zr����8�U�MO�� dZ�2�k\?�����_@��2���Ѵ낞��F��r�p1�[eBx�@�[����y�w`cLD�ws���{�OK���lf��/|� $�4Z�i��y-YמP��7�j̡�G|��U/C�^�R�j0���H7:ݥ8e�e�b?�������\�_O���^b�E��TLd��R&%�/ɡ�z��@I���Sc�m�Z�Q�%�Q�
���h�� ����X�@|�|�2H�T��`���j>�0�����l��F���׿���vh��4�U�LEv��5��}dԄnt	e��b��q�0��O:�{s�AK7:1#�X{4�u�$%���L|�_���j�]�]顛��OP*��1X}��jm�Ӡd�Z$�t?jQ�04�l�ّ3��)ڹ��χ{?%���/���G��H�gk�. R�X�\� �����Z@�5I�i<է�+Aţ@��h�z��	�a�=1D�Ã��]��l� �i��V����I9Չ��Ǐ����RI�+�;��-*+jJx]-���P�S�}IZ���x�7�+8�=WG#����c���$�v#}�$��kA�mA��jp�W�Ӫ��
M��J��'f��}���';��<��!�]�L����A��X�&��.Ɗԟ�W3�'@��MGkQKA���M��C�qD�c��5�go�;#}j�6�����˸���e#;�L0��
a�u����p��%t�f�h�[��b�7�MQ�H���@KH�{#~y����ek:��4��ެ�����w-Ǡ'�,�������I#$�&*�΃�'���`�<��a�^���|�n�}��N]�����GQS��Y�2������p�,`Ґ(�&d'0Y���*b����5�
�C�g��> <�<Ug�;�*P�2%��ҧlf��*Y����f���!���+oګ��SA�
��Fiţ� ��Z�U���L��C�=��M~�m�!�l���cp4l��l1^ � X.��]Ň����]�o�X�L������i��l���(�0�-9�\�q31ZJp�L�	�sǣ7��9��'�&���$�73�D2g�f`�;��G�A��r�%�ND'��k׺�gٛՎ�e="Ƕ�רձ5.��hH/��PC�u�)k]���w���+�iT�꽙F4������2L�
Ɨy�g�a��2%����z���:�M��%��rL��ӑ�I���6�=L�����i���T�a
���_�V���&�z�C��J���z��Y�~�.�D�����m�����8R�ͼXc���t�^�����Q�8��٦�A~��������ǭ��؞d�3�=L�J�yl�D��P�
t�~H�_�>_�==�.�O��xvm��n����4�G�D&�=��.�Ҷ�/9��3���pQ�e-S1����z�<��}�$�#)��M*v����s�r���2��"g���`�'�QR#x)]�b-�oJ��%;ZhK���^d�r$S�:�u$����Sʑ�1m<����X����d��T�F_�H�*�	Z&xޏ ��W��)��Sܠ��(F 
8E74g&���-ɓ��{��B% .���D�Q�uޠ��	9�D~�[/���:�+w�)�]��2H�LՑ�n \�o^� �`a�;���6�N;���Y*���q���_B�s�2��8��_o��2���B�pS���^��p�Ⓚ��1H�&���7Z�ɄӒ��RםL��B��^�r��ta�e���������C��&7o`����6�������=o�=�F�Y��qݮ��6Ι��W��= Xna]���Я
���1X7��dF��9D6j��~<fn֧���x��=���A����ƐY]��~F'7:��
�����,��7����1�������d�ַ��fQt7��#��{N�Uf��>x�,�C��&q�4��V��uO������2�N�Ó#�����޴�D�m��o�F���$���q��&��r'�^i� .�k���{���v�ǎ!�d��+!2�3HW2��aw=Kj��!��F�P��+U�FD�<�}"�XUI<N�� 6[bߢ�/��P,c��PS�k�݃�3C7ZĦ_�i-k���M����~u��俤���e��y����4. qp�^=I�5�B"�a�Sn����gl>\b`�yŁ˩r=%�㽵�w�㾟�AC�kZ@�kb�Z/��.�S�(3I�A�5���^����C�y���?\utxatޜ�Q'"@_ū[j�|k6ï�K�m���l�&��Y���.(�*d�)B�?W�o�{� �ŕ�ZO}��%p���:�K6�6>��t?������MD9�${f���܅���p���U�=��c��ϖ��ޅa��6+�W�˻���au���:�a����pq�O|���x,�'�4�B��ʶ�j,|�bt��lnr��k�����]D�b7�b��?	F*7ݨ=���$U�|��s~��	�`oT5Kx��C`��}�Jܩ��4�yޛ��gշ�����S�2hсZo�Y����`����-=b6�p,J���ݡ�L'a^\���'�ɷ��*i���bn3+	��C��&Y�������9k��tl �5eUJ�,��]�11�h��R�XȖ5	�d)r�\F'6�yh��C�po<�͈��!���6cC����w&�H��򚮟��Y|\d|llF������wJOsU��T碪�*lyp��K�z �s�(ܽû�����*����P�9��.����pRQ���g;1�j����w���]8���2�u�'�Z&md���HH�ع�
*-�Pg�-T�N�[���k�-��}���D�BU����_��R��֘���s��NI������I��)<5%X�$y�-<�|,�rh��a"�j� ���ϕ0�G�/H�"vM6X���x���Ja�j?�Y�������ϭ�����\,�ӊJ�
�Τ����=�I�x����h�q�]�ЫXF)��¼\u1�����b"����&�����s�(���%M
N"B7O�,�����Pb�.�"1��"L�r/!����-���1�w��h����Y�4E���xx�&��`�jӱ�?[�_���/ŅLN]b��#0��៊�߇���������~���m��?���}�?�d�����I�<EC�=�[�'� `��ܚi����_�_��·�,�i8��}�������� PK   J�X'(�5W �@ /   images/4737cce6-ef6b-4e79-82eb-dab57378d86e.png��?���?��*�N�Y�"<)�J�q)��+�9/9�ͩ*������i��"����ls�a�9nc���~=���O�].��?���t�^o�wL�=  ��߿� 80 �<t�w'�#ĕ�c��]}�C�O�!�������[� ?v�{Z���n���<�{q�>}��B�
n���O�;+@^�?�5D� ���~Y"}�~J٤��@\�,�m��g�;�o��]Q|z� EC�J���2q�D,�۬>�Xk���i�_TO�h������T,��@7A�}½���_ؓx[+��3<�������9�X��,v'�W�K���R��2���W���&��0� ��ِ���MA��+@]A�3JY�`���=Ɲ][h�Fq�M�p	@�3�Y���>j{~����;D�oy��s��-��y�����'���������߷��o���۾�-' �o�����������Y�w���9� ��2H*T8jfVtðKݠm�촿�h�X$��p�Y}���03a�H910�aUv�;�bg�"�gC��wf;21�m�1��m��K���0vTss���t�bbf쒻����|��F��C_���\7�.�2�%+���Q���}�Ȫ��dVO���7Kj-ڲ�v�S�o �>� 6{H��@��|��k̰���D���Y�>%QO�Kߚ��;9�ܠ��ܯ:�E��g��"�4TfIW����^�m"�ck6?[��;���qz��Z򧹤w��� :(z��P�F�:�G[\�'#�vg�#jKKʸ��Z���W`zb��+A�쫯1�\~(�J>�T%c،��&��ݐ�N8����_�h�l~��}�BU6�2���|!�`�u�OЭ]mz�V��"�����"��ձߪ\nC#�M��E�`�,��OV��H<���dP��)�����t�ӕ����E����O�.9a�q���:�bug���(�B�xg	������T_1c`T���Wcɟ��jܺɉs4�7k@$W,y��.�h��<^R�Wo�!����|(��/]�{o5Hn7�ǔA����4�//�蜿���%��6̋�)�J�6��7�a�/(N�˻@��wмiL�~�[�SLi�$S��q.�b7�_*-���j��Z]8Dj�'�^����cRe8��_�=+ZS�N����X[��MuF$���I/`b���=�nboZ�A�z�����n����42�����3��9��5�^CQriJ�>t�֖�q崽�j����֞EsV��,�(��>�u�w�8�$1�L�sd_�s�3R0Ոn���������r�bZ� ]߅�3�i�w�?��,oީ�����R�Tb��4)�@�{��u�GvލZ��GL���^>~ڥ�|u��,���Oٜ��W��Ij�̈L/|^7)��d�̰^��҈�	���y���	��v`�_o4�}��;[zoå�\B��fk�4N.������s����Ы^k��nH~�p��"�!gb��T\�{�O�L��t�K�Iw�����Rdl�d��B�oR���e�m����D�����h�qC�����Ҽ1.�*�>Q�>��c�8�
9�#��DVB���o3�mI+��5
mT� �hR�2��a�L&|Bn��^;���nM��}hq�W�΍��s��*Ʊm^A��xy�ڐ���ã�_u}Syk7q�	KeΜ���mC1*"Sw�&���(VT��-��>E��EW�t��ԫ�M�ce�.6{I�H]�sl���9�עQH3Y���KϦ��*��.Vj��g:rb$f�~��	m�'9���S�Z�Բ�(��2�s�,����_l���I綧:�J�B(ra�����l�.��ɬ�h�������H�v��/	��´"�8
�u�O��A��3V��3� {����|i!A��WNp�Ah��0�"�����yC�Pʾ���U���.���ه1�9IU�-�v�_��|�ɑTwƥ�0���۸��Rh��љ�±g�ckt9��OE��Uֻ}c��M46#5�2�����s���3�wNp�d���}-g�'�w ~��+�_{���UZ���\�m�XiI�7�r�'b����d������Z��'�t����5B�:Q������ti�-ܧӔ��0 ����!�ݎ��#G��ǧQ��5$�KO.�/��ԣ�P#�Ẅ���1z��]�C�>Z� �c���	��J-�ʺiZ2�xT�����@�>��Ӫ@��$�Gكg��on.���;y���Օ|p\W���E7�R���>9&��j����)�ѩ}5�$^xF��J��
�P/H�����a�w���ͪ)�q���Ie�G�
�dq�]��2�CBv�f��?"������U_I8�ڳ���4�R��� �}A�;-4S��j��:��t��<H93�O~|�A���M*�&�s�@����"jq_E/��1+�_x8���T�S"L#�I*_Џf���;��T�d�MSҦѩc���I��hj&�#�~��L����C`tk�� >`db�7�x�2CE� n@�Eq!�@�`�8W�׻'�w%��Z��<�������vw�>�,ͷYd��P��}�hy���qSǐ7-IXg����� ������R$g���l�^�|�j�6"�Mi�$,d�å��r���\�ۻ+~F�B��M#����͉l�����,d�B�k�G�^�ɂh���]���Z����q�Hx�C������ګ��f��nC�?#�d�<s)N�2U�RX�g�lWz=!.��H�^a�ח��@O2�,�����:�6���\g~�	ix?��z���\b���6��.rRU�u��Y�t"s����ya�4�����H5O�)`m'��x�e���n��fF���%ڪ�������(�{�7���}�L󻠫�)
䘱��9J d徵ΦtNr:)�=�S��xBN�[�9��S���
B�L�6�٭���'3@fKe�0����?��_�1V��L�����j�!��#�b6�>!��9�i��������XO��c����/�~З���eb�nj�.�������ey�F.���_���+���H�8�-!~.��%�C������9]6lt1ьh��-��B�D�݇;u�\d��]��C`JN�Q������AY�X��q���S�Ry��֑=���$ ����#�o����T���F�T"��9������i̦r�5�uٱ�}7�}T*ВM�q�Șy����ـ����!\�S^��&�)p�´E�<�_8)�3�i��m���8\��{i18W�u�Ɓ�M�5M5/f�Y�a��~wr���;�s �Ҙ%��|��REټ�#9�W��㼪�?3+�2��z�d��#�-'�"^��������Ra�}Ϯ�j�>�w�hI���lB7����;�V��/$wv��=�>rRK�
s�3�	�宮�œE��,��k��x|����,�w&$�]�W2Z�׵dD���ywEwN��w�DX�aN)��F �*Tca��m�.�Y������]��I��$�}���=¬ _,�F����s��Yj�W�n�>R��LMϋW���=��MYP�B�|ٜp
�I&�I�z����039pp4b��2]o<��d�`�؞Тg~n~�����C�����j�Um�<��pk��;I-��͈ȹϱ���."��/�o,}�X��-���z��;��M��sQ�zl����T���I���m�by�hz��kqv�����<���e���%�0�'�^��BN��� ���5���@,�v��n.C����hf��Х���	a]a���Iޟ	e,EO9�b�`��)#b�]���7
f�.���}Fl�H))t�)2�.]���9櫻v1W��m)D�2��[dow �Yx|�vw>��^�>f_��]�ߙ^��s7>�va�'s�ŝ��{1�1�4�ЏuW*���$��L]�>J�@�~A|��)ז
׵��A�~�[�\� ��?)'5�̗�{4{h`!�1��^����m�	�{��AeX}1"�Š/�����[ooA)����}r��Ŝ�}p�i&A]�P�Ik�F�F�`k�����RXx�T���X�i�X���]�^д��k�1���s�����3�5�u%�T��u+B����a�V�x�m|*^�^�g%�_��K���vֽ_��aR������h�����y~$6 @����k��{�~�%^�xb�o�����V2c�����9�6M+tc̦,3���M�ww9����.���m+n̥��B`=Y��bĶN�[$��o��%s/���a-\HqJ���sS���(Xg��	q�F`.e�x�������@�"wܬB�m��|�.�Bv-�_,���~�z(�_���b�������č�Kގ-��:��'�C��P�J��D;�Y�ON��)}/@o�xQX��t5ؔ�P0��u�Y-8;�EN8�*�F������n�>��ó	��x��ƌ��srZ
uHX*WJ��:z6���K�g��ɵ#�V�ZI��喱
1
�ea�e��j���c���!߮ ��Q�����AD��!�����_ת
�G��R7�6��O��,����L>�i����^d)O�s.ډ��MJo�����gh�U���;"G��bi<��$*�2�E�N��ԤS��}��@��`Rv��%͑nR����9��chU-�5���{GWt�-�$'�=��"����ǜ�k=��Ij�ɢ� ��J�ވ�y�~��IY�[	��/2��R!|��4a��?�����+éO��x���Z�G��_^^ܣ��M� O;�r�Ơ�$�X��c�{ �N��M흌Ɋwhi����<��s��7��1o��~�����'��S����!���:���ئ��'�6�7YM�!�
 �F��F
��4���o��"x�Y3�"U�r����i�݉�oOن"u�c7��m�����H���*�A]SN��<�1vh�����)�=1�Tb�������������Y����v�֮�m�/��ɀk�������m����FП�c>+{		��UjV;/��sx�<�8v�V�
��d���/�Gl�*Z�C�|wがQT""�ioTMء�^��Q�;<<Ί������X���s�~�ǜ*y�~'7��N�d����Awm\��D��+周�e�ɉ��P�z��C�k�I���\U�V�Lu�~5$�K#Ex(�g�%.s�o����S���\�F�{|�cv�����n�^\�69Q᳦�54s�����1ƣ�9v�o�ho�ՔL��Ȕ��|TYZKl��Kd��J�WC�%wY����c<��ؐQ��;6�����o@GK�[ܩ��߉Lr��h�(J�!usD3�����s��?8~#yg��t���~��Z�̫49$��`��KŅ]X~�O��q���.�<L�V���,��ǹ�J�.�-���cvn|���������ƞD�����>W�E�YQ	�ח��y@�ƪ��D�����p^N.�z1Sbu���*���İ�U��:�K4��h�ac>���m�۟0�W���ZbGޯ �_�ym�#qÉ����X#�=wnb������e��M/���v	?h9�N�!���j�i���=�7_��cby�#7�5�џz�g�gy�95�dw��'����CJ�S�/ic�Ãe�� �]���8y0 б;ڄ��S���t��A�icK��O���V�*9]��曖0��q³��;uY��3f/�1!o ��V\�:�z�^S$���)x��Q����
�UL������|J��Y�����/��sVY5G����i�^��*sL�J�q+�f�\«�X�P�v�6D֯G*���!kI���\�Nl�SŖ�zΦ+�_%0�~����R7�&#�7�y�oN��t�n�=tp�x7[�N�C���h�j����F��Iק?�)ğ3b#��܁����W4����O���d�Tս~�2�s�g�p�7f��˱IY���f�^�N~�݃����./*�:44�)T���#�/�<�/y�'ܰԢ�� _y���i��#.�n�^�9;�F,{ȩ4�=�����.{I)������r�4��(CY���v��_�<(���/s���'F� ��ޟ?N�~��=8w���r�z����I׈�'X�6u�~�,%m|���sҜ�y;{w�X`��O_��bҁ��VY��>t�
��skŨ�f��tR�T�e����|���`���49��9���2�^�~�l���ˍՋ���ٷ�q����%/���w��R�~��Ϲ�z�T/mp�@��w�5j�~�y�%9���H�O�f���Q��و�P��T>r�7�����>0x��8�:?����r�&4Z}lI(��$6I��$��2р�|4�;��'mt6����'2�op��+Msg)��jՂ M|����	 ,|OS�1R8!@8�-/y�ߺt�7�'���-����I�;�.�OK�C�a�jw`R���vSM�DH�$ԑ'�o�vQ	�CN<�_��h�A{��A��XU�BsG�B��bHY�9�rh��.�����.G�b}��)�M����S�x.y��^1���*y���3�D�ڜ��9ިj��f۟g��鬻%�,�1 F�|��Xp�b�u����s�2���� t�������hB��8+�좀����y%�Z���.󿑀=�^�Cb��0�#"ě͋W	9���OT����� ݗR�{��")J1&�T]j�J�aþ�l�)?�?����V�i�ɦ�y<����'D�*�<a�d4���GAD����r�w��-Th(:�"����"���)�uu�ʁ��[��fM೔ӥ0����]?52��-�� x�u���������}��5_ͷ�hx(�����q��;�
�Q�\��	h%ۤ�(��m�����3՝���T���s������H��+��Nq��M����ˣ	m���G���(jE�gy;���7���'`�� D8z��)��cw*C*�5]Y0�|��r��-�9$��Ϙn�i�.2�
Q)��uv�(���\�Gh�紨l���o뀦�)4)�\�o]�r�@U�Nb��eZkr�(�{������!�?1|�{P���d������)���kdF���6.�H�lZ�����W	�����	9x��. ŴD���?�봀��T%א�,ƆX�����ZC��4R��}冑���ť5,��Su:97!
B�hA-nQSיMAs�ugjlO���:h>�<�*���à��C~c�X�錄�X���O��X/���_]�L�3U|���|R����Dt��Ӱ� ��g���������˲m-���f�u_�=�i�ꋖ.���
Q�	+B����s��J��~�n�-���;��r�p�m;1�'��D;3��jEt.n�� �����/_��_�������3'���(���EK��$��í,�����@��z���fQ0�_��>���?��0*��<"z�� <[�'Q��^h��w�c�~(�L�����\T��{����~�a��N�f�Z�2DO�֗�RXJ���N4�R6x��"�e��Զь_+�9�,/���}����E�Ǽ��m?�n�q�ո=��!�a�}��6 ��=���fч'�M��j+�P+O�j/)4�|��`�4��U�!C�����6�C���ôl��LCO�h��]������Ԝ4����6Zo��L�b"K,�/�k����Ł���
3���_d5t���fD�(��6q� �+�`���ol�^U����~�>O &�/y�ϵ�w�V�u�y�t�nο�ؖs�Mg�T^�Rӌ�NR�����BBdiZ��Ρ�$�q׳�[M�'���C�ۦg�����Aҏ �ҋܗZ����K,�*y�f�syM]�
\������R{(�{U�ȅ��Ë+B�R��*=�ۀ�O�A��'�(q�z'z,3��!u�Q&Xp����c�����$��s��n¾t��O?�_Ij��p���`�v�j8���1#�bWL�}�oK�7L*:.O �o�׬������$t����7$L{y�=86}�v�bb[�RK�KK���+����];��sssWh �����;
�Zv�Q[_��_Nj7����R[���7:p�*�#	�I�k��&��]S^��2���:%��9��[��J��H2�^�iVONd��1����u٣�FB6}NU�Fmp�!YKTmbQ�1T,����iX���%*�Ol�_W9�an'S��A�4�P)��7��Zx�1O;3�G+4ޠ�?�ɹ��H9��s�1��2~jkl{Z95j\�O)���p{qj���
]
Ny^��d��*����z,��9���?��~����{�Wݥc����8#���Ps��՚߽&:q �jwz<R ��Y�qW������˷]q]gQ	���9&O ��o6�5R��|���Q۩k�/>E�e_��'2'��}΢�<��8S���7�f_�,��sW�Lb�F�ȥ�z��MHc�#�:"=� �����q1�����X`@�&hǩe�V�Qҽ�钷j�K"�fI/���� O����hT5T����>�9��^O
e��r��K )ó�ьMqz�EP�v� G� S3�(�q#�̞+U���9
��}j[Om�7��Y�(3�v�{��ot^��;9*�q��C���G��������ĕ=B�z)?e6,��X�Z����JS�[I�M(�`�J�ɭ��^����DU6II���0����w���_�c.:��Q� ��L�"пbc���ȑ5�w��>�1�X�*����c�ڃ���WEed����ࣗ3NO(=�F+��\q�bV�d�~܃�e���RѠyc��H��L��V��P�^�wi^#�����m��̻~�@!G��PO�٢�N��{�~6yY*?)P<V�Ut�va|*a-v�S��a�
;m��i��3x���}�n3CX�Y.mX}�Zoc��/kd��Z�|8��􇴯�s	M;w��?�W~�����������Ww�v��%����Ň���|
?Q{miz���'�Ow�o�y!6�t^�|6_���lߧr=���B�����9o?��g�8ROդ9M��I����Q���g� 3M�֏p��� ���A���s�7�m�0m��L�0T��CA?�rp�|�d����)iTg�Ͻ�	���r@��슢��SMXN��<B#,>Q�ˆKp��\�L�-K���G��d�1�$���q���ieaj% ��]j�o�-�Q[���K ���
�9^$�h��2ΌF��������_O;t�6������� ����	�>�*����6~pD�܇`�`�=��ƕƅ��28�J�p�!G� CI�������s��ǐ�zY�?�<n
�A���:�z���|,_��Ӽ-��#�@���>��@�m��o�.:rH�G=F_]���p:g돐�+x##|�a�^˖�X6W�
nFo'o���[9�ƭa�u1�vWX~ڰ��  �k]	���r����mz�79_����N�k�j�	w�� #mTO��ZȜLH��(N|V�Q��dr�����9�~�����AaxM%-��[B~t�A��y<l�P!����Ƀxл?n�  ��yc��!,�!��ȩ�N�����I��_���RW>g�8�*��K	=���>�8�㈱�i5Gٟ�dv.�n�2�Ȟ*��zO�G���\`��W�K!��[6m����,��K�v`���]Qȣ'd�yq)G*��.��.Łjұ���A�)X������'bku'�"�c�2؝
�o@����[$���Ƭ�7�-�+���.s���"<�u�����XI~�v�mI�1Dn
,��^���^H�{��]Q�D� �����
$�{���݅�K\ V����BqRp���i���B��5�	�s�!F`+�{]��	�7�(�{4���H��7���Xb�����xf̽�yfο^��OAV
H�ʁ�a���P�0]�z*�=��2�""�}}�8�Z��㴑J퐐�E*���e*�֟}aegg'�{�.~����V�ڿH����+��7S�,��5s��@S'U��L��ը�0ݸ���o�?����$�
4Ʋ���С�'hz:c�����C���Y�RifT�b�v�Ȧú�~"��<�ӊ��b=�D��B6�1Q��Ŏ4{��I��	�����E��>>���M�M��V� �W�\��O}�r����/�>(�RW{�3�����x+*!141�e�����7fR���5�^��kuL\\xlͮ�LN R͗|��N9\X�`�#µ	���Ek��THQi��=)�8�6_9y7��f��r�>�g#����?g��3;��i<ox�ܮ�������XH�����cu��H�������� �-��_��}�j0�q k߲L����9�\\��^��?G�6�zL@`(�%uV$C�>z�Q:���Ij�=A��DƆ���"3EJ\p^]g���^_�'5A_�Uu"�-Жg�·�@�;��>��<$s+y�	t������sg2Uй8���=F�m���|#��ǎ��rV���My��|�i/��	@�����^��,l;�A0_�Ryg��v@ߡ~��u~��8�u�b��%���/�}�.6c���{X\]�X�K�����U��\Ͽ����?�)f�1�����^��NR� qE��G�����<Xg����].���N=R���!ja��o*�e�R*L��������[�rj�=�P�[TT�)x�|?Ԑ�^�?D���(��Sg`�ǉ?��j� ��ʨ�!���[m��m��_��׻!�O��ǧg�C=��3�(��o�m��l��
�I&&�H�#�i<t���'��Ŵ�0	�W��c"�$H!.��<v��|��0v��6!�����������.�E��}o����g`Y��i5غ+�G��0�e{��?X��Բe銃��a	����x#gA8�%��0)��#�dO����S �p>&�恄���	�-0c>n~��� �[Ӂx��7���&߅��Co�m��,���#�2��)2�ou����l�qy�m�Ѕ���O�<�-��Β���+�ˌ ��EQ�#4x}�|E>ux�D�s�'em��F���:���*��l~�Kl���P��(����ɪOOW�>*�<�(��'#�/xIQ?߈"��G+9�_�}=�j���-����
^�����ȼ6��f�bx1,�J:�(��[�S���h��X���Ƚ�F�_��7Cu�	��̧�����e�}^�����JjRUb#�'��� =�Xz�v�,)�Bح��s7{&�W�C�}*Z��aצ��2$j��ޱ7�E���� �����p_H�v]�ZcN� 7`d���!z�{����8�޷@s����k�?Y������������|�ʤ�o�|�?u�W^8���O4����3�o9_��h��,%��j~A��s�G4YF�,;���[�_d�7P���
�.����PRR��N��Ø��/_��j�?HB{���BK���!��:%iQk�W�^w��.f�ܲ�Bim^ck�{�?v��*dD��|Hn�A{rkg��TÀ3�"&
�S�3oV�4�4�`�XX����ٶ�Q,��C$��8mg���$���؍!� P�7q
.�eK}�񣖢��$	$(��'}0|�7�����{��l�o1�q����j��#�;}��"PT1�)ͱR d���A�f�N�ɰK�=�G����Ğ�P�5"�:��=YS\]=�^5Ը��˕c�!��b0Z��*¤��7�)u�Ch�<j^Jr�-��C���T7�����Kd�(��Z룇�������ۿϩ���զ�g�\�ޭ�%��g8͊��#�M|U����&p?�wu���CZSէ�,Ｖ8�.~�r�i� �дy��эO��?���R[*�=�	�/�l�]F���m����z�`���ʶ
p���5�fW9������'������*���ڍ��~�0Z"�A������JG����Ɲ�rj�ֶ�|�/y�Jiٚ��*�0�2i���
tS�92*�Zz���ohŴ`mxI�,�=J���mQ%+d��L�^��#
��N.��.w&80ŲyU��ɘ�G4��W�@�e�h�T�?�O3�WN�;W=X�|�.���)_hX��,7w�H۰�!%����H�tC���ߢџ��ME�q��S��gK,�4n�K��v�D�[IcJ'��={e߳Ί���Y���r2�0�|����E�?Q�,|h�l������G<��SF�+�D`x��	�*�&�0���4��+Ф#���h��D/{�x�	o��>4S�w�{�<��v6������7=����&<*.*�}*�Φ��20RL6_�x�Wɇ�_��.bP�uV�Fj͸�k�`�SJ�g����[}}�f[����t�U�������r�2�v���O/��
`桩��'	7��S�h�J�GD)�L���K�e��g�1%|w�mN��u0��l�i�y
�V���t<~e�˛�
n/�vJBRC�I$R�o$`19�^]���o�T4��d~x}��ώӻ�< @c& ����%�BXt(:��7�T%/k�2k�a	��@��J�
�]���!���AK�Ű����\�B[z�!��o
WUSU(������zT�TИ��� ;���UL�"�jb2,��ШQ0k�\���)�m�e?��6�a��I��B����ꋇ�R���J�}��НL�����+��ywd^>l�	��~?��uJ	Ainv�ܝ�.2� �x��t�t�uɍ!oւY�!�<�
�X���PB���*�K�V��"���^m�i���'y udȢ�0L%�Q�^����Ⱨ�6[��عǨռ8��3|�3c��zN4:�
�ߘ=`��h�D��܆tSW��{Wc�s�!Ý���ȗ� *����h�I=鬋���dK�%��~��{ı��%��www������(��z��n�&J}���Fh��l]p��uʕ�w�Ԟ��T&I�����?��v=�}�iYf�>xB���se��To�/Y��Z��ļ�dMZ1�-��p;Y�?�A�1�k�I^n�ɕ�vW=�[��*P��wX#:An����.�t�Ʋ�<7cE���wynv6�_�E�FZw������?�e�p�p݂Ka��)S:�gF�r��ᓘp{R��=�6��u?w����.���i?G�{��{N��)�����FM�������_���\�Ǝ4�Dߔ*�:~e&�0M�K,i��y�m�du���só���>Z=$}�lKy�ְ��N��6p���6�w���J[037�#��s�civ���(qK�U�A�ST�.����*X$�P)�7o�{��n�eh6OĮW趒�+ӌ��oT?����U+�nL�~���$I�Q��鷀����;�s�?���\��lY�49xk�W��---[�`���U�-c�8��F���3>�tujsR���ր��Xy)�	��Ϡ=G��ո cy�Q�שd����R<o��ϽR#=�����t����[�Gm5��VVZ�ɗ�Y��P��;���`j�����;���(��g���&�h�3NM-s{�f-,\P3r�LQYi??)˦	N<z�P��tg D����
!f+��fR�O����)��pc��EK�k�Xf��&��1Fx��Hoↆ�V�4�@ �G{�2|_�n��ȥ#K�&��+ޮ"�ޮ���R�����Z:O�ڂ4�Z�:�[��roI������{�n��v�`r��m�����PR��vwX	�@y\���9�k�4

"���l�ձ���ּ�6`�K��-����
S�U8�2A�9�7e�sH�q5���p��@J�Y?� J�F��e�իW����`F���S?H��t���$�ݾ�ߴ�:0��ѵ��C�nD���ɐ�kw�����o�q���J�@�_*�����U̱+���Z�A���4\�K�(U�"��=hg�%a<��>M��@Q%���U��'�$�XϮN:'�hΏ��>�2�kg����}�e`3B?��]���Z�b�����GWA-�U����BK^)
m�z�~��)�2f-"���x��<N��	��|}}Kȡ<&:Dg�y=�
\�����q�����~l�}�Q�V�^o�a�j��� ]���jJIf����f��������pf�17�pV���F4����w��CPڹf��:�HJ3A��`s2%���X;5���h���C�vGs���FDR���@�֗^E�g�
W��w���4X;[.��wp�&���lc]����a�YF���,����XҌF��Dť�p@��}�ۢ�dd6��M��I2k�~ސ�B%��3B��4\�.�]e���
\~_�XF:�P��#����YV�)z�%��k�a޼�U�ߣ�04z9n�wG+���+�����%���rؗ|O�?�r����Pl}�})�BC�zZJ˺�q�R�dg�Zw������c+�R��|���f/���U��C�yn�`Q���Kz��@��H�MH�OQ����3�P�{j�X�������b�:��߃���nR=:8ܴ�2-F�����Ԩ�W�"�E�"��]�/!U�y/�\���U}����'�u�X�Z�\�|@Y�vh-~�_�x���
0�-|
��qJ�o���E�w$Q��i����R�ȯu��M�_Y�ʭ6ɽ;Oge�۶�B��RQM�5SʴvN�ph���!��vm���_c;�/C��j������8�G`�<
�򱃧ԑd�6iL��,uYb��B'��\�VZ����T�@x83�b�jkj>� ,�a��~Vc�f�7/�a[�WK�|�����V���=������TC��iÏ#G�ի�"#�q�+���9��C*����>��}@�J����!S�%7b�̾2A��S�];�Py�~��|V �gY�~�Q�S-��� ܢ���ȑ�{�4}޲�I����Qr�Қ�?L�9����̀
�%�;�e,�_|�N�2X��߻ #���6��pP��}(B��4@�������h�VeS���h����z'�i^��`��v�O����*�H��Kaas_RC��SZ[�9��.���Y��:wR��T_�L��E[��C� ��A�X���@4�a�
���`n���U�6�=O�=-1W?����î��^��6=
f�حK����-..?�i�eA�;�"�7(�ÊA�*��Wx��� 5��8;�t���{�qur�9-}�q�_ݧ��N	ol:*~k�􇰡-|�"�ţ���� ؃W�Y���rj���j e8�o�˧_s�Q�ي����n��+l�	�n�ƹb�F������'k��Ƥ�W�s:$�I��'��l`�`U�Vvl1��6�^��"$R��az���CXicꈦ�j|/{��#x?1�4��l%Y�eETh�eʳ�,��n
�y������uK�H`h���cjf����l�#�9X��J0�3;����KS�3��Ōeo���e�k-g(g�,@Qd�c6C��.��0Wp���P8X
^ t�5� Q�'?_��q��q��]p/��N~���}�y���z3k�AB��e�gw9Ws�|��g`aI��MtD�m�fj�� 3n�F��:�Q�m�`��5s���t�cu�'��?���q-|��W����͝����VI4fH�$�������St{Rl.GC�o�(p�QP0���4�Ԥ�w/u�YPūqovӑ�-��ձ�N�X;0TJ��X���0Ib>�`�a:�d�����-�N�����L���H�fM�����9�/J3�a��`^�I�=�N��y��P�����;�i�Z��2jӱ�H�O������`-�S�؆<�Q<�z'��q�~�~�wƏךT�֡�O��K-r��e���3�z]�� 㼈�O�ѩ/0�O���ơ���U�]J��!���ٗ�N�U�!A�?F�+Qs��=��j�8q�/���	~1�v��l��QZ;�[�Sc��L~�# �>�LK,\�0����A��TIH4H��&V�����S�3!���j@�W�����kN������G�/V_�?iK"���[��غ���}m;��c�c�)� 7}��ф�kRhƏ��%���@E��M�cZB��b�A�j#������-����j�
:ʚ�YL��O�$���ǖ�j�ۅw�mvH9�٥��v���%�}����*y���)*��r�q��[|��"�8���ݏa���h��s�	}���N�Ci�{�]�Z3�K5��mz���L���d*��]���ׂw;�������#Fd�7����g��,�=.<���+ok�j
ߴV;�`S�dV�V�6�.��z�x��[����`������*�n櫶L��>����<�����/濎j���RX�
Y�Ⱦ�w���m�
kZ㦻�C�ST��9���H���K�k���e��Q����N�<�}
Y$����S]��J?�NO��t�PԷL)[�Y��L����1��qM���8)��%R��))"�"���0:�Q�K@0�FKI�1F7�a0ꋯ���x���������{��~�$��"]im��H]#Rj�~���^��mk�2L�I3���q�G�T�L��=��CD����hM*��>_[>(`����Ŋ��HCOc<��F�7��Wu�Wq9h)IGj��:�Y�)�!Ă�rS���MvV�~��Q��tM�%�=W�Rg�����������5�V�x}�{XMܞ���B�z\2æj`���=�;%����IxV�[@5+��Kj�K? �\/8����I��!z�1���M������}�=Ǝ=����bjS͋샺mD�T������38��P���/뻳qR^�k��L���tS��p'��P���/� �޹�7b�~oi�"��/'&\���0 Ǖ�G���%���շ����ʗX�^j4�4`���ĻV��f��ӇWJ&��z@���1�G�1Q��t!�Vg��>sV�����k�D;Ƕ���]�MYh{N��)_q��6|r�E(w	�k�'%�*���v����N:��\�dLg�g�O��>ϗYLQ-�V��%�œ��8��e�͢���.���{n���;eʻt���m�= j*�cfw��SH氛�几�����.-ޔ\Ej�"M�Z}�R,��5��nsX�$V�$˷4����yz*PO��L�X-��{-�&�x_e�QB�@�ȇ�f	��m���;�h'�:�)�X��=�=R��|��gH���C���7��/�F)u�2M?cbZti�\»��m���e����ˀ�I��ȫ�|� -�6��׾�R =����1��ߜ3v��mB�ކ���\���3�i�Fm��n��=��7"� ����8��y>�Ɓ��Y4��t*�{x��8�����c�g����4��U�"��j��iT��s6�R�8
�q]�	��U-�.A�����5���C�r���=�}dI��zP�������U�͍�`�ۦY}-�j�G��7rO6�{plνl�}y�� �:)X��sr-�r-A*� T�rf<� ����!k��U�-� �>��I�G$8��s7�)�ڎ�+vi�g�w��Q�����Q?�R�?�;�Î��4�*;/�>�}zt�n{�%�tySFEBok˗�l�e
d�^aI���y����(��Aӯ]�b߷��2�>�`���7�?9�OӶ��l+�Z5X���خ��m7}�S�TMX�v]7�,[���b�ٯ�w�R��)�����n����ڟ�#*�,
IIМz�����U�$q:u��,�F�Ļ b��5I�'��:��!���v���4�3\ϷZ\m�I�Ȭ���I��q\�]���U|�r�Lw��J�?9T�!~��a�;�׉��	Nr&{Df�d���.��v;!��{�	=�f63�c�P��(�kDy3,��G�1���m�d��)�j�X�̛h7�?`B�[��&��.zze��~˷%!Yf򋷐i�8 C�{���U�E��K�7����W'��]�^lPFz����q��d���H�+�A9ی�w�5Y�-��]n�P��m<��W��-#L����2F7��#s�o"�+ey�x0Q��7i ������m	g����״�8�6�ac�؅��yn��S������7�V�n#�$Gv��|���s�.Ur�3�9��QUԀm����T�z���z�"��(cN���,�.6�yߧ�+��z��9γ��N����w�T�qZ̊��)�j��Cۡ�̯@���*s q�
f�7"�~=�6�O[��˻�^�{��*������@$l�~[m=�L�/�Z��M��}_	��_��4'o�P^	��`� &��(+Y�6��Mf�D�y?%O�n�ch�_t�@�-�
�%�;_=u�X�%��b�7F����?�ݖ�O�a���F�2D���\k�O��ϕ�k��^��y��{X�x�r�b��|d_�mM�9���G^5H\+���\/7]\�4�f�~ ,��e�3{n&���*���j4�ֹ*i��)�;�Q�c��ۘ緋��_]��C�8W�st����}���A:b-�|i[s��Y�ޟ��B6DL{K�}^Q�.	��r�����+;�;@���=�����4�L�m��D����M���.�Oze�y� c����6격3�)3���z(;�'''�J1<�<����bX!��||�&�[҆&�#h.?7W*�����g�pX��B�w?T�8��rrdI��X�̨������W�+�q�,IO�"�(��������T�_��1��2y?���7撑N;u�:���u�p,r)���)AP~�_f*H'���zUWLw"ڤ�� A�w�; �^��Ҿ�j/�J�z'���r��1���4ei4`_�*O�����LN�?-��ѷ��Iy&Y���#P�� C>c�6��I$����/#�Yȟy/���!���Y����R�|n�B!ϲ���k�0�l��R�9�ِ�{��X�s���m�iJ���̏����Cn5�9�*����)��y��Y���T�FoY0��Ol�A�!����ا���a���>����Ͱ�:\�" ��~����w��=����cYx�Z�1�M�H�6�ߵ6�����c\�.��HF��/���?�{mVz�Yfg�{�z����(�mZr!�y>�(QǼ��L���1+$_O@��p2h�@��.g�CS���{�w�H�!>aT�.<z�'��%Zuq���J;kx"���b�XeH8>���@�5��3ļ�/ۜ+��G��ݻvxw�c���:���阷&'{nfO��t�(e�����n�u֘IQ���y��z ����^�RCuu>_�I����;��[��I�A�5x��y/�ֆa�e�?�����<g�_�R c1u�U<ţ|t~��ɘ#�*,�u>�˗�a�}��s�n3�2tINǅ��!�k�m���M�I����F��-R��с��W�u��D��u���F�������-��xMR.��YUP��>�S&.����o�L� �oW�a�뵬
��0�z��E�m���4��3�xG�ti�|*N�e/5�Iǅ�����6�1���T�����Nh�uq�\b�|���Ad�5t����:b��itd�^�y�3���e�aT�2��B�o��w��.���ר�c3pBd\85��&��U���"�2!q$�� ����u�_�}!$E��`s�~ Yu;����*����g3���lU����x�HY�7���1#q��{�^��Y����חQH)��uV��!�&�6�lZ��M���&��2M����+G����c��H�與fn�Pa��C����u^�_z9�]��Q�W�I�Ǵ�E��>�ң���3&Gh\
�H_o�6;|�_�0�uq��y�%+��O�ڢ38R5�s��jcndM��-l�,zCP6�VF��.���e�`f���p9�Z,����>��vk
�YЍ'�J������f�J�Ϛa��ڑA�7�2�h��K��z__ΐo�e3��xL�h�|�[RRBc�5ӧx��ڕqQ�S==��y����CgO��M�m�H��MB�k�6���s��'�D�L,Dj�e�W�иԠ��9N����~5C_�����7/]�e�0�5:�����I����3��%�_�s��%��pq�z����w
~ʛ�M.*�1d$+�lRvx�Ej�C��U�Ł��^�s� g�&+]��Q����Q�R�%�т�ҭ$6��QB���x�dVG��5����^Wb�ti��oy},����. Kf#C���^��g�č�N�;-���5i���s27G�����y_�^�{���k��߁���eQ;Nz8�S	.R���$ᤍ�Żv�=n�L0��-��;����ׅ��g�!�a��J��^ ����	!v���Yl��0/}HV$i�`��8�y:ZKЅ?�q�!�5����{��� ��:�h]��1�f�������u�[L���9�]0yF�ޛ_��YP�@�-��S�(�&�v��E�3bݖ���~@��nm /�Z�N5 �b}��ثS�3i9�r�}~��ڗ����xjF�V�ϻ��N��SuEmaO���RvP���ݖTS S;,�^�H>heۜ|L�<��~5�(�7�>�G���Ʀ���h���P8Wya���	��I��;���YL@0"�j)\�6�+mn.j,��� ��0{G	��H�����/�EÃ� �l�?�[�k���������4�^)�V�"� Z��L4�����I�̬�s�3���9���d��)��>3fz���"��ȇ���4���&��)b�%�S�yp��%;#Z���V#���k��Z@�Q;'|x�s2qkV`=�ǪU�Q��!-N�7�S)�2&Zk�w��1O�C��#ɻ���=���4k;͏���o9�$�:j;r�N��q��$��'��i*h׻��O��(i(:Ư~~2"��v2�`r�C�~�_FKyܿI\"�y��v�+}&c	�ҋ�>WJ�-���S�#�������
S��9oS��{'�����(5s|0(�S���i���{�K|@H$2_�sz8��ڨ��D:�����w�xٛh;����i����Ww���"���M�ڹO��;��&��;���)U��E�2�Βl�&:z0����z�K��lu-�!�#m�ô�z�#��]�o�Y}]OWS�8��kK��2<9��穹��,8s&�6}TЬ8��W�p����Wk~
�wQ��N=��8o��oI0�g�
Z���E��>�rs���
��P��s��"��=�P6��zZ���c0f52�@5�pJX�@����	Lh�N�Ɍ���-�s�>�8�"P1��������� ��7Mƻ��
�� ?��5<���΅��NY�F��l�MP�̭y��5��y
vx�7Kɂ��s˒�,�?���y�i�Y��b'�Y��>��и
���<��y��{V�w�:ۥ�x8Y�^)�K���dn[��z- D^Jj#g�J���"`1\h|���U�&�U���n�b�c�3��V�K���%�P�mv�ٹ��|�v�tZ�c��HXR���%l�W{Wo��4u#&C�0D0� SL^��/;��-;���E���\%�vĨ���lD������f����6�7�*�q�i������ў��D"q{e���lB� .���3B��nd.�!yNQo+�6�N� �b���ڇʭ�X�Z	@Ri�E�Oz�'m��h��5�2�Eb���sT�I$\����C�_��9���3r�{�Ag�������!JH$>�=�c� ǚ��.�q��EH���K�Ѽ�vv�������s��"c[���E0cx��<=�������-�Yi]�/D��f��S�[����gIjO	0�$��)�+�iî����m�n�U�3C��f�� q]�U��l������S��g[!���كW��5>¦���b��-���U�=O�|��Xy)i�+�st�٦�D[��{�{!���I㠣m��|䳑�Y��sS+!1�z;���c���ov��I�B+��z�~������G��:eu�A�1���/93i�^|��>Y��d����� ����.:�����N�=9�Y�ď��`���m��ϔR�:D?���}
�0�\�r�/��'�x�[�����VK�&�/߃Bo�>`�8�*��0|N����P�4�m~Ox��j���D�M��dKhS%�6��
�O:�K��D��_Q�����A+�:IDHasE(��p5�f�f���8���}�r��)��'����ŕvAn:���"a+>��ig��4,\ml�]�W�J�{�0r�����%������ϟ���á�S�<�5�+�s��٦�H�8��QT�����3��^X%�XE'�r*�B���t�h�7O�e������:�SL��|��d�b�e�������D���#�Y�R��pM�������7F��_ɅDoE��1HT?)l�� �~�l����-̢��Ha`w�IC핡��39k?�tn�Ok|���<�V�O��ҩ���{��qW2$Ș$������0�Ձݒ�,<Tԝa5en/U%�P+9�m��Wdf9zӞ��T�� �ۣ)3�.z.f���cgc0(L�mFy������w��z\�oU�蚹*[&�7Җd�v�,/� 	��M���%��^ p|u��a����Bj���9$�]ԤQ�9iS�.�M��H%�}�p<S�rᑝ�\��G����9�%�E��%nխ� c68� ��n�����N��&���$o���U�C��ڣ�/¨���*"�W�ߴ�J��]�6��쾛�}�&�$�*�Ϲ�yk45�f����lx&qv�
)��%~��zG�h���H�G�ܢQ�9ܡYq��޳i��N�g�րm��Ja_���V,��.ز�6P@���7=���T��^��ɾ��런�ݝ�.��:G럏��
��*ͯ?�f۔����z������ŞLz�*�sP�Z�ZD��*����+���S�!�n�HIoFZ�}%��t����w �x֒�r�/��3Q���݈��l��ɠ�'p�'��a#/���x�x#m1�ZHz�����k�7y��w���Pk��ů���Zo�S4O�����(����b���o�R�vTq�"�d=�;��Mu�.5,T����O?Z��i٩_fǗ)h3���A����J�d��������F���B6	���PH���֌)�q����%C����?s
V%<M	�R�4M�	(�L�2R�W�E8����Np��>�6�|ʖ�b�W��P�$�nb���bVD?�5����W�<�#��N�G�҂���R�=�VFF��A�{!>�V��	�x�3Pϴ�zv?�z����l��bY�e��e���3r��@��*��]ϤM��w>�Ƃ]��NSS�5;y������G9W�G]�ȸ��=����(KWAA��Ӆ�;�iaq,�@�rL#�7yS�|�����۹�� �!����M�����$;��Ë�E���Lo�������_�f�av~�[w��4.���4��U��,Z���'r"�"�څ�8�d/���+y�ȩ6a�l�|�<b���a���+?��Tv���p�W�1�2b������.�li��6,�󋜄LU��@g�Kk�=���h�]z4�}&3�� A�FC�.�"�oV�aȽ�#�,�ܽ}j����]h�E�>�(��>��J뜜[{�L| �c��>@=CV̹��Lc��|6���_�c����I���lǧ�u�2g���b4�"�Ԙ<�1>���a
���cC@�d���XL�GO�7�+2Wg�%�n��c� �Ii�dN�.B�F�_5EO�L)- �9Ae�LP�W~k<Rd��PU��:���	�W�[&���
���'�x�?Ak~�������A�7~"ծI@!�V�s��@�9��y�s־���ҫ������;��� ��Q�V
[��8/A�5o>M�V6�2�bڐ]���x	��n������O���ގ>���Z����M����T2H�|�ۑv��L�8���i�y������ylz$`:���	D��/�mя\k��~6Y&�A��c�}&!jQ�r,�뙴�H��rز�V�����h[�N���	?�_���Q��EȑH��Ǥ�p	�Z�4��A��>�tc9R�g��맛����*��n{:�-���*�?,������� 8����<Y룢���(���"i�5nQ�7��)�n�2���>]�@�O�\������Ԃ�����踳><�ʴ6�JUԗ-.�)v�`/'�[���'w�&��fd��~�<�^]6��4;|��^fJ�>���Y�')�33�����b���<)�U���~ŷ9Q��93ɗ�y+��+6�_��̾�1Q��6~��_]����U��2�m:C<���r�|8h�*��0�7�%0���w��(���0���Ű*���{ &\'��Z3�����ui��+��!]�&R�E먀�ϸbg����ՉpK���*����@���ŀj������I����.�#�����,�ǯl�=��϶��zc��B6��0	X��;��o��yt�i�;����b\h(:�I���>�K�Up����[��n�LJBY�?kq@������|�On[����A��"��,�-1J2%;*&�0�rY!_rs>�.hG��Ӄh�w�Y��.����vo���3j#XM�x����12�/�oX=�Q5�ߙfO�'�@tk���}�)r��#�铟u�{Jm�0�����l�v&��q%@j�/�˚��*�mL��Zu��E|y�Q�9�(	�Se�tK�~-.y��&s��kf�5���Ռ�'�uJA_�\�����˺��O�9C�Rs�*��|��qئm)h�on��h0�zz�y�d��\w�sl���}7?��F��� �r�H�ix/�rd0D��=/�\�Z?�!h����v(2xL0�з��H��~E�~����p�NiΫ��2�����%Y�ۚm���^�&<�C�ACC�������/��N��Ϗ:d�$�nI�5�_��[�������!011�k,�gAfI���+L�i44������@2ᓍ'�O�Gjk��G�Jn�u��|�q�Glb��b���)�7ɥh��W�=�f`�:;+����37/�t�M�{���XK�M��H��[�7W��Wi"�m��[�A�X����WI,���O�H����6������;���⃚$A���?=
Ꝯ��\0?w�Rڄ��~�ԉBƑ��wXE�J�{_ס������N��y���6J�E�`a4>Ʒ�e��?:�)�҄�� �R'�4�g:�TA9�|*�^ �r��Ls���zK�j��	 ))���3�g��^�(Aw�L���؟R�۶ʵh�l�+Y����H�T"���Ѽ�� �Js{�\�#ONN�Y0l��qԵ��ǭo���Z2�AR�,e�ǮH'��T5����������م�X�Y������Ϙ��s]�WX�W�pc7t�>���N�"�׫u��X�h����/���G�E0�K�骈��;Y��c�T�Nn߼uk��S_��<ޓ����n0``��|idC�i�Ѵ.�?��9�̷c\\_e���e*�������*�P�ޤ���}O1�Â9�����%�y����»��@s��J)H3�({]�r�qBD;��Y/e91
>�Կ�n���q�|ً������&�_�8E�ggh0�u�߭��
�R�+q^��E���w��L��p*n��+�<]��!×�&��B}�����M\�Aں/2c�f�m!Wl��Ni1�>���c�vT�z�o\*'��Os�(�����IK�8Xl=�h�\�Q��β�W��]��+��![�Y�W�D���4].��R�]����U���l�V��=va�GT��&�	��C���T�]���kpaƠ�-�U�V������B�υST�&	T��O�O�L��"@`�s�fx��F�l��U�
i�4IJyi&*n*�D������M��FKV��μk�Y�,u���33,�)آ�'<"�¨~�c���T ���M��V��'�?y���g��-�h�!e�^����SƏy�8b�������;z��D�oF5{�<v݁���fˢ�w��=��;���X���?4Uh�N"���{�Uvzf�[G�sR��Z����Q�,���B?��D~�iJ7�mɥ�x�ѯCt���ă��re�Ptu�b���)�ǅ�~���SƁ�:MQ���������젡�z�Pp�tt�|rڟ�m��\�Y����wл:_��:)��xF��!����Nx�g>BN,{��C�л�L���J�0��)�H��	�[՞��~��4�١�9T��Q^[�d�Y��j|�|8��n�� ��E �?G��<7,b��c܄dM�gLOw��u���ӆ��ג�f	���Gj��g��һ��Ţ�]�(��]���5��TQ���F'�caC< �΄@+�{�I97��H��ޠ�>k�ڠ�56g���XN&�^��ˁ���Q��x���rR0{���Ѥـ{ò=��>b#�@-ǆ	�z ��K��=��\���������:�(�,۠�������'aE���ܼ�:���]dß�� �k���'b�/�x\@���
�֬ճ�������,��O%8X�	�z�����W��&Y1��Y�����î�H+�����^�8���]wQ���;�(��/��4{<�Z�J൙5���H�]]HQD+��1�T缷ک����!��g,0wW�T��v��o^�ރ�v8?�0��5O���`��������z'���1k6)|��-����������i��I��2"{�5�V�_�ޫ�bYȨ7���6�M�2��m�l���<�pRٯ�-�f�#�D����@����k%{�\K��n�N��7����힥IjR1�}�6�at�j��V�����P��N��`w��t���P�ʿ�Ʌ����n�f�B�����bg�O���_�J�t%��[���R���x�ػ�q�����}_tM.��jh2K���ėe���}6��xp��L�q7�xЭ�f�x�#����&`oD�ۚ���Y]n�F�&1Sā_Z:��`���Y!���n�ǭ!�Y��'����Jׇ�R��Ҽ��ge���f7L"�.u���$������}������I��m�k��� ś��)v�����A��!� Tmɕ��ə�����+��,ꏓ�����%e}e�zo)�������Juvg py(����+�QVsS�d@`�g��io"i#��}(�XPk�;�U"t{��R���W_m(�ݽ����v�eх'm�b� t��qҜ�k�N(�K�t �`��=|�@~����J%ʁl+�Wj%�+�(�~��<o�6s��Nˑ�3 ��t��~�S	_-Z`ɻ��"��Y|ڄ���#�=���-���@����C�C�9�����2�qsȟh���o̾G�H׽V�n�� �5����V��H9..ߎ.����@�)z�?z��`5���ɡ��z麟#�$9�7��dJ���쓊���S�n�	�\H����D���Q��9�6L�jR�ν0o���s�es�8���{�7�Ǽ-H�"�@����c2ls�q��<���̣�C�y֚�.�Z� w��~�:V�iB�k�+�ř	��u����wq_�_��ij�R��d��6�_�q���b`W轿�Wb��}ŧ|��hm���H~QY4��Q��҄p?|�����W��m��<@�+�>v%_99�Z��uҘ�+2g�B�ā֨7x������p[s���2msю�,}����dQ�{��Z�`�E��Ϗ<���T�`����s�wR/Zeھ��1���]D�5D����=��B�(-���[��Y��=�����Gr����;Y��K,_9�C��[q��PQ��ܶɐZ0��q_޳�1�$����󛃡~�	����
�J"%���9D,G��Jǃo�?8hIHb��0�ha�s�&}?���}�n��Qz4�����G�]�X�*��@:�9���]��ځ�����iv���'�j����'���1P�d����	�K�+AUI��7�����}�t��5'0�r�%��7�'���M��5�^�8�l!���5,@?���������޲��f���f"4m��nŮ��VZ�
�R��K�uI��Q�bd�I��ݻٜ,�F�3�\��e��0x[L
����l@+�M'@%�����Sg��6X�Y41��'���h��s�O�����pL�@B+�\� ��z������ۍ4ȥ���������%ϴE�5{�'֯:��Ka�^0Y���/_&�a�n���aެc�~X� ���ʗV8!���R|o�״_+�.�7!�a�w���P��b�_B�*COK֬-��5��y�K�@ɑ�/L SEoJsY?��'B�r|ʔ�MB����՛%�?�<R��[Y��)���!+B�tk�2\)���~�1�r�����G���&_��[�7�n��]���
���%��s1b��A:е{�J���'��#���0�6>���#+Õ��Y��e^�AiZ)i��Q�A7�wTbc#ˁ�),ݭ^��6��@������jm�(!-=}_S�b��Y�����ϧyS�e�x#Ekང��Ox�X�繿���=uD��-��d�o�Zg/�Ĕ��Mu���mut�����e�潆�l*� ���N��ȵV�4<�����7i����b�$?u�i����c���Ƨ(���,x�6Yi*ΨL��Nȿ���%���b��rt�/��v�I}��b��fM��1Dv��J�~^����U8c�KtR�Nq޾���&8/Wu��W�~�/Q,I
�O�M�(ǎ��>�I����?=���h>�E�'ᩡ+"\����c�Բ����[�����U�՞����w�_���H��I�8�X�E_�r����eܟ@5���EÚ���w�>trAt&&&TTT�ד<����;'/eo����clp� �����U|��r�^�`�bo/���r��
����fX�{��B�Eg�\��QRQK�^�Q%����(A�[���v`߬ѓ�}�/�:�Z�M'�\�jX�-ʺ1׉Z�aP�	I������dZ�_�bēy�P�&����+o͓��`���2`�����*�jy�@/#��*����	���_���Fq��)72$�(����L��$h�h���*�}!.Z��4;�� g�tz���/=��b�ł��n(r��H��bC��i�k{�����xؗ$��Ό�����Zz1[RR�/�Ӊ����N��j<w?�76�����m}O�(iM�$c�4lv��xa:99]��u�nmm��T�Z�w������PL�	�ϕq�5gI�_7���m�}���ƴW���e��ܕ=��K���c����Cw�,�aq| ߧ�`���2�y��+��i�䜈t��t���t�&�� �~ɱ�Lw���I�'�(q�{-0�Ν�d����oWI��B��p��w�6GֆB~�<9�Ώ�C!�X��o�DҢ4��B�s������X�wAHC��{�v���+t�>��,Új���r&uglܺw']���G����\}��ި=!�&/� D>A���ߧJi�*U�a���/�8�D�ar�ÿA	_��K�<ل�P���K��
X�yNN������l�靏�+U�t���U]w���\�^*o�¿a��/z0�'8�Z%Қ-�%��y��2�߽�]-�ekC��Ȣ��ȗ��!�!$97���gg�H�e5E
_��tϵ�~���]f�-R������`��O7��e�ɥ�4�T���9�ס<�����Ofv���e>�fs���>�5�10o!��{��\1I�&ݸ�a�3�3����3M�I�������y}��*���4x��h��bg�5��y���!�鋼�P�����1*��ôP�z2Cզ�JԦ��$~l�䉳�k��z��s�M5P`9�����;���U��n,+��w��k?'%�����e�6��5�eS����i}�;���������-��B�@�-:�***��I�P�I�2�<�28��r�>F��M]�w.��k��Ƥ���+�'�T�Dh��l����UT�s��.�z�i�b�ҕZ�����9�;�:��\�N_|5>�AV�Qύ�?�{\�q�o��f��UD@bY�-͟v4=re�U��p����?��c-n`���A�[�/�7�l����DԮ��KJW�A�U����L�� =��U�����/�Uf�M�$�q���'�X�;!��u�.}���;g�.����Aŷ�:{�N�L�7�1�=�4�*��h��m�x7�,IÚ���7x��(_��O0�=;�xѴ���#��m���LV��Օ�_f�؇���o�!l�3�ey����ϴ<6��p�[�G����=������dct���%�vҩ]ME~�l�x��d&"H��6��f/�\�0O��"H�r��(����oN���qa;�Fe3�����فi3zΨS�Cam�c�[o;#�$)�;oK���{�rk� �E��B�_��.]%#�Ր����op�b������w���`F�XUz,d�d=Y�MA��U9,Y��
�i*����[��
?nE٣����l�&
Hgt�X���dzr?���YT�}5��$�,�jK�q� �X�0����9�յ
ʊ﵍�z��#,8������[�}A��M2��Rx������a����h��8�����t4+(-�N�q�TkQ6���t'I�(��V��u�o�۟@����	�����1���%IIII�38Jc:����6?��}������S��=�$��}���>% ��|{a��OK�ge�
�!ڃ��Q�:�pw�(��+�����6��6"�)��(�/��;�ے��urPn����D��)�Dn�����b��z��B�Sb�VDe2?u~�+���J����!����$\"\�Q���ř�ր^��j�B����Ʈ���ꃜb<�ޠ���XK�}E���Jc?�cW�}�$��#E�=��]ߛ�n��K�MK�"�	��nO�E6E�'���
���h�Oag��s��穤T�>�y�ƒ��JCkJH>�����$䭇�"��Ի��Yn�>�.�r�/8�V'
����;����3��[�t���w&F��[�?�/��e�öb.�ޤ�[��>�[�-�
� ���I��.���	M�,B-6_^o���L�#���kЙ$!#9oiE}��'.��-��g�$* P���m�z��  ���/�!~���ET��M�:������F�� �ae�@B�ٻn�/�Zo�ԏ����cL�M��Z�;M��P�/;LS�@�F�*q&N۫��S��s�߄��b�M�6��7�\_mG��?}���.ķ<��̌;b{�c|"E���%���1��	?w��k3���@:��}��v��[ca���rK���1Vq�3R�D3V!��y|8v_��q�pm(R��;�!'��_i�h�`Ӊ��u��6��!p���VVB|�
e�v"�\�Pw��>Q_U�4ɖ�����4#�����ᓖq��
&8��Y��4Uz�p	^�����U��*<�u�᜚e;t����C����
�����j�$�~�F��T*�+Z�֮�J��ܷ�N�o� N�ԏ��eY^�]�Ԛ~�ؘR���`ȜS5�/����FXklf�S�������Ӏ��Ml�/�Ы��>=��oMT��l����r�s6�Hh�(Y_�թ����"�?�5�h]m�?���\�Z����o�Ŗ�����*�lU���ϐ�W������,��� ��4��.7��)�)�1/�ƠUtQ�
����C*�#���=%�K�P�'G�,��/a�M�Y ����lj�~�l9&�l��MV��&5:�N�ѡ=_�}$��Nﴣ1���_��7��Y�F�x���|O�J��:�k;�R���������`;����66���>���`7˝O(^{��<�ۓ�����U�௓��*�B�^�q��9�����N����I73��u ��s���|"���NM�c�ۨN����/~�P����f6��ÛR�LC��A�Y��*����G�A�s�f�����e�G�䌱�h:�?����9�5c���5g���%�W_$d��N$c#2��h�
�DX\���;�>�rĚ>A��Uq����:���
�頝|� J����Paf�����'���*�*��c �ٜ�	�`>���f�F��憟Љ�����g��·J�����@��瞥�l���Y��dț�D�;�d	ݼ{���� ����o\��4^[�S���?Try--�4>�����ƵFAmm���{F�?��F�vvw˼2a/3eھ���'��.­?$�Ey�r��±�x2�_�;�]��Ѝ�/L�h�~��[�����f�z�>f0:ϩ��L�]���my^�a�s�,vg��}=�"±���A)&����#�jP���uv���Ez�p�Y���'��:[s/���.=�p�E��=
�q SRhQp38�3�I�͑SZ�q���%�9�h�Xô4�'��up*^�R=��"��r҄P��^W��h{�e/�F�b���Ks��*�o#�HRE�s{o7N=��~ؖ���I��	���‛-��������8QkzN��٭	��d6tz^v&�`ܹ��e~p@�X[1gX׿= �����ޞ���?����oq^�%f���V�լ�W�߿������]���������S���1��Qm���8�)�R�w
����wEw/�)��]�C�νg�/��/�w��=��y�0��1Z���u,������a3X�����:٨��O�^k��솒��y�����<�>���&�d�A�m�C5�nOş������J��T�B��CP�_-f�CvZ��'Ũ���I.[|P�Ķ1v�����d��#�#bC<� ��t�	ۓ*�<^�Z���M�ԌZ�����g�$檌'{����{�`�����D��,�k�?�F]M�eFw�.d'DC�I����@O?̠RG:+�T�
)���h��|�w9��}����h��u�umr����>�CJP��J[F���[}����Vp~��l�{��ٶ-�����]�!��Z�������_Ҧ5����/f�m|÷�u�� ��Q����A χzs�|��z�*�O�ը��,7R�����D�[М�`���\^�D�Ed�Zzѭ|����/}�����������i�8X,��>t٪Ǘ����4��%���m���	���Ĉ�]�8�$6G:xLXn�xPE[�J���b����Y�|2����Ss�Z#6���ݩ$�+ڕ%LW j]�0k���S�~-{����'f8�mE�f;UDw;�:�[��F��`3�N_$\3�@���Jwu����2��y0dc���p?�����,//�Ɗ��2��Ӂ?��l��5�[�뿔u���]f�T�, �OA��>���v�d��&@w��O1�C������WU�w2wJ�Jc�gTy�<gưEf��g���%��=T1�{ԑN��\,�9��B6r�Ǟ���q��ݷ�5�_���(1�V��W<E��ր�k8!c-a�h�	�oa��0R�nK��=�%>�M�w�f�lV��S�Y�]9�f�#�`����{�ScW��(��+֗vq'���у_c�\@^����h��"]2:16���
�F.�'1yr�HZ��;:�^��VOT-!O��JY�{��\�Q-XB��/6���	9�����m��[�6����<?Y����r���-m��Ym;.#����Ûy��f�|rjJ��C3���F��;<?�I&}1���)|ZT�	����X&����VA��=#b�W#�Q�;D�4�k�ċO�R�P䲼�:�6::�ҙ���`�&��bm�ɇ���VvW��v�7�Lȴ^´+��f�ؾ��C��]���G3�"��n�Z_�>�uu~�: �M�$�o�=ɆP-�ʙ�C��j�Q�C�Y��5;0��6�� �h�ƈƇ���xH
�t�����D��� �.1s�H/ �\~ρ�L�03KGܵō��xiGƦ3kU(��w�#wf�s�u}��\�)Z_$0ͬ�Ӿ��\"a�8�����mxv�̿�b���x�ҍ�Ņ�������k+���^��Uo��7�9��_E� ��`�������/��8;c#�>i�ֽAt��^�U�E���i����l	��6��=#Fsd$>�RS,�_I��gV��h��m͢]�G,1���z�!���l����lܮ���9�3�~��fn���z|�����&I��X�F��^3�Q�.��I���N�|R�c9=�i����V',�@� ����PG������n��g@��y�K��u�����8��z;3g3�����-�\��0����׹�k�;":��cv���b�D�Dp��(;-D�
l��]�0��ҰG��9�S��xƌ���r�ۭ&V )�c� ?)��U󲽜�IEbO�*���6v��������7_���������J�}��{��Q$<�2~�

�kO��зv�r�� �]���/A�Zo���{U<w2����=���E�@������%�Yh�����z�����B�x0�3�J'���:&~�ݥ؎c�������+�@z�p��f�Pn/��l���%fr��	����l��}���0;q���Ϛ4�e�Cx���Lc�LB4C5��c1Dv-�5��j#R2~�m���ɡ����?�;�4ֿ$�k��O�h��s�Y�����:Z�}���'�uGO��>��x���jmsh-G�]#��uz�+v����sO��ylw�ܨ���u=X�v{�5�B����H�������|qc;��?���tg=-dm����� �WPzŞ�{+[۾��o�K��U���	�"�*	�B�w�xb�����Ȱ�ȭb�Ö\q1'����b��9���Kو��XTn�@	�]n�w�L�;�Yg��q��1-&���ӗ���]��p^�S��kw�Bn�u:��\����F��]&Jt���׷���qWVr��ul$�u�d%��sI����Qb~kw㘗�Q�:��L�'�Pg�=��i@Z2�v�O�����ǏbL��	��m����w1SM�A�����G�ߩ�Z{|j	�p��"pm�|�}t���I��G3x}�C�V�T��QV�Ħ&��NX����
���������WB?|낕̎�E�J�v�Ը�M�3G�̓r���,}�j̽�a�Y+������uFGGk������wܶ�n<ݮ�93��l������]��f���kLGGw>�r'����v��#�/����:"7�K6g3�(l�6��s���OZQS�"*H/�c�Rk�nP�|�1�XK�-|Z�O�� �9X�Er�i/.����m`�~����7�|��y�el�I!�����A��웋�2�����cy�-�r(�o6��8a�Zқ��՚�M��ԛ#����Kc�},L�bs�ab�y8D��ƕ�r��%��r#���>�L���ݩ���gPt���s#��gvBpi�t��r,\z?����K�}�ݎ��Tk�DgH�ߠ
�2���ʫ�fbN�½����P���Ԯ���������mB���v���e2|��`���s�*���ƞZ���)`_�j��A�J=�Hʱ��&��ˣz��ëX����WNN�k�f=�%���B�=�`����k�����:�?����1~������쏡x����ZL+�-F䙗�c�=:��d��d)��^��sdt�Y���Q��]����ٲ�ak^O��G�Tp�PP;6���o>��@PB��C~��=���U>[C4��p-�+Щ���kl��|��$���~g�%��~�d�T�#��1hD����)�t�s��m@��*IY�9���\����cF��jS�7�]F^�tur��b��KS/����~b���c<�b���)2?ÿ�5�`0�M���zYR<H施6}���*�9>��ǲ���(v<��"�P�S�润k��C!�v�����FJv*2�"�R�^Tajcm��S�+l�U��}�/.z�jQ�#�_�M�+S��b�]�߰y����y�8���6ⵇ�hq��Nq{�tJ�>˗o���U+�e7��/2׷ �)d
�^W>�e���+ͼ�玦�l��S���<h��⯬���B7By�n���K�!]/�NV���t������@
T�frIgl�3�����>�Y3���!*&�Y��[���?��cf]�06�����9u�pf������� �Z�ԃ�^�Y8���1K
e>A����Lx&!�7�b5�E��KGh^.�ƍp<�{7յ�@+)�6tϲZ�=��h��"B�Y������qoX��WOk��щ ��!A�=D.X/����¬����3��!��z�Dwr��+w%��rqg�`�������-8��oQ��ɤἝ�>�`W4A���e��x�q��S�O�MT�LA�iY�� ji������Zy9���:%�Z�f+���w���������u�DSItEm��$���j��6����
$�rk
d�6�N{f˵'gg�\���1��8/)�/�V�W�%F6~�\X����rN�-]���b	褗��A�Tb�}PEM�]��A����g`X�Y5<�nCC�&���A�C�WA��V}?�z���%H�m��%$"���X��U����\A���|Ꜯ#B̒v�|Wzʠ޳�e��^S�� t�#�U��٧9R[��[��0D6�e�>d&��a�ha|�x\X�x��n��sb,��7��ǆs>;�U����)���+fC`\��V��B③a+~��=J<;�����p�u�6�F����E�>�����6�d-��� �α}���˴��4{	��y�)�)���IݼQ��B�l���ej��w��.M�6��ZS�΃n7AK��[Tv�@��2����ȶx\�|kp��tC�>x�6��Lɻ�kΨ�=�]"���v���"�5�
��#�T֤�5��HuW�ˆp�(����J��������B#`Ygҿ�y6,q����r=�j��M�b���w\F��ǋb1\�/V.:[vE��3.�*��*Cqy�F/�m""Y�����MY�����
�f�!
�y�Xu��,��ˋ>�V�o��z�=�	9~H������a�h��$Ѣ��p]�k�|�6��v���}ؒ��?a��J�`8x�c>L(���Ɯ�.
��9ݹ|���S=���5wM�U�5���PY���ExV(��/=����~�m�n1�$h/��0���I�c����B�c����.�ZZ���1'T~�3�*�5��V/�u�>fp��K��) �a�m��a�ƙ�&ۛ�68�a�`�ה��M����� �E�*`PC�ɒZh~���;)���`mԥ���H�\���qn%��4�>��y��S ��t�<
r��=�Bba9�?s�t�)����EO�0+>�F+�����n�����|�u��4��3a�௥�q>�1��c����Iݦ�>����F렙���lF�nn�F@�^�)v(
���T1��sv����i�����2=QGG�(�ޜ`ͯ�bg8�D //?_m���}!�|y�?=��薎[_���;������Ӓ8�m�8��!2!�d=f|T[s��VR?k�eӓ[1:��'�i�xqs�8��(8��7�\����F�\���L!iNO�=�s���VH�s�2��~�U�������(,�8:�݂�z�SO�s@a�����/b�e��~��tˣ��mi�i�K� ���,h��r�4���CTe���W���1�ќ���-:���4|�#��㳌�zZ��ŀ��#�0�_�dG�j�?EݼR��ѓ�����y�b�ع�"�h0�L�b����a|2Sr��|:y���>��������`��*����1�_�0Q�w����tކ���_g����P�ڱ�1e�X�&z�r����X��MS�]g�nW�曝�1W���� ��j��w�_��.�-###WۭuX���L����wd�d)��q�WZ���/���n!%ǣ�77��k���'����Sē@!���1��'j��j���+a`��;j�瞾�P��q�6����"��Q���r�Iq<K^��0uw��n ��
>1�Y�NvY1�R"�,�Y��zu�@S'3��
�/ܼ:�x�~V��J��[ƞR?�$[3�1|�@��Q}�{�Q��;M����V-�iq�����ؑ<mU�, �DHxcܻ�I���ϕ��ޗ?�Tvo�k�Q7O𡒟WO&7F�\�A�̳*4�j�ko�a���2�\��ۯy�b���t$h���Z3�=�sV1�x���f�x*i�[E\�ϲ�M@�;�CW��Ӻ��z���B� KΣ���_�Ɇi�P�I�o%�;pR?�]�5R�^z�uT��Bjj��k>�2���O��d7_�� Uo�$��Ap�
��	�\�v���Ԋ�Z���X��[�r����imKM�W�rMBY
����L��}�8��QX�U+�v��=j~��C�!68�ĸ�������vY§��^�������)���/>v�A2W(�,����>�tA�iv_����AxR�U&opL?;�p��M�5!K-_�Dk�8]����zr�b��G]�<�r�6��19.���~��q $c��FOE��peQa���iC�`[��N�>��}���n|��A�F�,\��of�����ӆWU������G��	�,�f�k��[���n����-���(E����
S^�-�
9�����B.��f��������Ɉ-�Y2]^T�rvd9^9�D�1�}�v�#\��;�$V�>;����j;���I�^�O=�� ��cc
�WE"���_hj�}��Jk��t�k�q���C���wGR$�6��?v\�n䄒�)**��\�	�2� �4�i��!/�ȿ?�Ujc�j2#�������Q�_�hj��W��'1T�d�;����A����y��y�PS]Y�\ۑ����+zk�+��+����R��|C����Ib���~�����(�Bw�Xyj�BTհ��ş�D����͒/B�!�E�C=��^q@��J�Œ?'��VYқjxEQa�F��7?J*��_%�ɉԆ��y�z#o�-������7���(��a�`��g���Rz+��W����l}5����u���0�E��{e{sȋ733I�),��e�kb1����A�U�����/�}�����@%�>%�c^6�bT������b��>�Vi��%���hRx"Щ
�Z�����q�}�x��)��v Y���I>���'d��S�X�pg(�8��u����~^�n�)33���?�6���rr�5~X"�U����K/;�7=�HX:|Q�(���U���qBN�:���w�+�RdWX�3?��'�Z���ua�?� X����Q�7=
.�hP�tH��E��nK|��� �H�
Y�Kq�&y�����^y���~����ѫ��A�A������
?<>(���m�c3)������
�'NzPMa)"¢���n$m9�/¯����}cm��4h���G���[�r!��~nN�[�a�͡cS��g��;��I!AZ��W�w�6B�950;��\��;�=ŝ۱r�z��~����y�xo���)�ԆQW�7X��N5�%t��HZBlؕu�+��\�<e�!��VY<8�{�+�5��ܙh�q�x���K^��Am��F(E_W�h��^���&�@����ci_�s�I����/��F,燅3͛{zɮf_��x����a�2 ��T�$8\�R's+�;;K�^���	l%�-> �U�;�j���0PxU��p�(Ѱ����7u��$�k���k�R���}�bB�L��������O&�sx%����R�^�b�#��(��x�{L�k����/�>�BN�[��w�z�'kvWB�+x���Бm&�z�L�,���<�hI#����ŋ��c9���
Z��c'V���oS�93b� �B�ho�hٵ2�4+`"�<%�V��B��P�M�C^��B�{��6�ЦE9<��X*���/v> ���A�3�|�YKm!�J�
y�o0�'�95=`�����}n��PL�d����/���2�'ÒN��sٻ�bn~�p�5o�ג8z�\��� �EQ!U��Q��K��]F��O����f����3��G�	����� [y��g�_?/��xu���x�wJ�R�z�?I�)���UhRps,e�Rc�S��)1u�8Bmĸ�ټ����Ä�&m�nOs�&R9�C�hQ�&�>a��v���_M���ry��{��.x`iw��ls�w��W�|���ؙT���{.p4�.�[�����s�'c�����Ly�'�8�{]=tT�b5�k��l�n��)��G�xŴ��a���8k6�]���cz]�o�h)���v�Dz[oTVD�j��5Q(�-8�o�ں$��)Eˢ�턎������&\@�Gqa�/a*�N�#Z8��c��]���ʩ��Nz&���)���K�.�z������� �����1�RQQA�+��1*�����gR����A���;����ۭ~�g��a���3��{p��B��+�y#���BK/Y��ͥQ��p��"{���!5��0�2�4|4$,�-�Mâp�|Sp���(�Y2�>Uk��P��]�ݝ�%�_I�qL�c����R�w-�2��?0��o����W'*J�Z��cM`�H�(�
>otlm�V���[$�$uM��T*���ě��$�՚���n�����[1b��F��&c���d���oȄf�7��ʦ�x�;:�EI��ѓ�j�Ӽ&e#�7}�<���wg�Wh���;k%�ύٝ�=vw��3K�h�k�81<r��0�\('�Gɻ�Ab��Ko�3a�9�r�P;Iu�9�BT���#j�V;��B�S"�k��uL�}&O��~�?��s�&_o�5��m$�&��hr��v���b�8pMu5�+����|<���?�JD���75e�ե7��y/95�ʙ����ֻ<���}��в���bC�_՟��g�\���#�o�&&9rKgHj�qo#Ҡ;`��c�0��Z�T�����D���,"��ē��>�g+���n�	��QՇ���BDwS�R��p�H�> �����v#�{����[/ªKO��<&ˢ��:��p*Vy�k]V�~��Q�`��3�U&M����j�0�v��9��$b�8q�`��X2�6lL��FsU_t�Z�R[U�g�8�Q�	0PQ����P=~kR�[���+#�N���OY_�z�f�=WQ���6ml<K���ey�����K����D:Y���è+><O��h��~W��%����>f3���\���k7�4T����>����a�E�ٱ,���gB������.�-��]��X���'%��I,������q��c�|���{�$�7\o���]�j��ɤO�� �4:�ǆ_��.�=�%O`Y[Qs�J��J���攕����AB�L0�
H��Mа�4�T�G�W��С!EcK�,<� ������N�y���oZF��9��IRqµ���c$A�E����^Bg��b�U|�ZpNI���}�Ksr��j�P���5gn"����_s�Y���}Q��1��D&�gm�gjI�}���ؕA�zsE�Xѕ_`N����8m2�g$?@w%��X��Mvdg=�w�lKQg�� ��%9��C?7_���I��-qJ�C�Xj�~;'O��/�W�n�O��l�5�C��D=dEA�k�l�v�����E�B{���H�\�?~�*���"���n^�Nb����6���.����z��+���5h�o�����W=ł�JD�ՎGdff��lQ�>P���'t����B_SJrKE0��}Q%��^^�T�5�5u�W�UrC�������p̢0>슏|Hߏ��^�����q���Ý���Xn �݂��%��ZF.���.�=�wR��[�<k�^Y��=��[���^k��ph�2�{[�8Wo�q�K��fl��P9�Ԩ<S����U]ƫV���@��!�8�ĘE<d��w(s|�/�;x�d���n��U٦>�T!���R�lƁ�q_V�l/��qTB���O6�ؽ��L�nU�^p�?�u��	�LZ�\n��P���yY����J�9��$#[N{�i���<�� uE�$�PeL��ӆ�}"򞅤�.9�g�ڸ��Y7�$\��n��g'��yB����B�b=�0Wa%3���	E{�b����_#�[1"�G"0&����s�,�c�g�	/C��X���&���y�&�D�{�V�_�2{��_�VlR���}3�C�P�s+�za�6�	�G{��V7]:^�4��#Å��D��{5� �ʄ'T_bHqB�����h��#.k��JY�����������������?|ĢT�q�Y�Y��{�Y�̬�T�.����*�g'#�Ã�`)ʳ�9�P&hw�%�����}�L6�w��]�ID����Ҡ���ZVғ�*�/��r�ݞ�s��T��E��#��;L�4p����50k�إ������!C�dQ^�a�?� ��S��f��6xX��$�sz���ɭ��)9H���>&�fTK��h޼$K����;27�m?���s�Jִ�d3�`��E�W@&�^�A�8;b��$�I�������~��Fxµ�_��c�;��8*O�K������Я"�p��UH�=~�l�U���K5!�q�>S�v���jpN�I���,ڊ��]�՜l�n<�ϻ�Ӎj(=�9]�p)l)���\i"��Տ��-�H��w��`���ZgC�_:X��Cu��L��!^"4џ�/U�Ju3��˵�Zwq6�c׌��?���,n�3Q:!��t�)<?#鷥W{Z��+9@���M���<���_ް�?5��i~_�W̏�?����q���H��8�n�k��(+8�
�V!<�ŵv��3{�$�+���ր�v}���$�x��]�����1��J%��>�HL �լ�^�0�E:]����Vp�--X�����4=�,�?��֮�y��{��~;S�K�N��`��ER��wz�(Bcm�O��D�]��]�ZJ�8[�������4y �sq�M���|��Ō���o����(�b����L_�H��{Pn�~�W|Q���.;�B���"�E<���4�=��w2e�*@�`�0�'{�!�3�t��ki/�'z�N���?�)���&|d��A���ܾ�L��8%Q0ti����5�5N3'r� �Lf�Q�`������L����R�_��$���y�E�����?Ʉ���\�J��O���"�Eíp�ȵ;b�|�U�	t�Շ�hw�!ֆ�׶�o㥗�B#� �p*ڌ��{����)�Q�{1Pu����R���9I��q=�g�3��4C�ckVh�2����2���C�i]�����?rn�|�3a޸����͕e�e�	lcdg���i9b��f:���I!SP����~�ӞB�vc�kYz+k+���z�>>>����@!���xe���4B;D�"6T�E�N�U2���U��C��<�{e�l֩J�h|v��g�L�~E겿���>>$�T�)��y��u�l[�<��f����^�"�~���]��:N8�3��r�_�^E0�v����d����ѣyHVh���e�8I�b|tkݨY��j���gϪ��*R��0�"]t�;G�E�#�>U<��|c���;77��{�L���(��7�,�]�Jf�?7�;�M	��w�;BGr�3m��1v�.ܽyL��9k>ܠ�(����O1����f����]�d�C�xg��� ��扠ѕҪV7�����Z��'�����5� �i�~��/�������v�	�+7�T~��&G(z�YJ���"���y�嘀�Sl-x�c��T��l����&>ׇ`�t���n`���eZȎ~������ D�ү s5���L9y��8���5�̔E��߃��+9�Zo$2Ђ�%��u�$���
�3�ӟ�����ۡ��d��VRD-)8Ṵ[F�᢭��ߏ�
�k������v�,��L1����:�z2���5Va�f�8lF�J1	����d�[��MSq
�y�z6�x؆��*�{�_6�}���Ղܡd<�u	[.@�;���c��x���ƍ�dY�|�������)���ћ�Z���-)��,7�#*j��j�d��8ݢ��g9MD�[�mK�VO�� 3�ls�~hx�o���I��m٩Vț	<x���q-��2p�$��!��W���B2�cO��������?���j��&�}�a�:���f"nkg���*�'3�/�E�t���I���p���̀�����~vv*�Y;����|l������	!ږ$k5�;@��(,[��14����J������:�(�M�)G�#�АV�B���8���	oE���y�\����g�Sq"j|JG�	�@3RYo�:�g	fEUeO�)OW�ʃkʱ�DS��Њ�����Ӑ�GG �%WER>���^/�pK��h�LWfY�e�%���?�b����-}���A�a�����zAe�h����! 6��ݍ`s�s��Ƕ�̦�����n�Y��p^<�B��'6�:7yt�)α�GGq��}ٶf��z���fg�*��!%����X��/:̾�R���̢��f�t0��r�V�����&�I�:����z�dN�0.>&_g���O{)��c�Ip�l�ަ�B�1T��R9~���8:�'T��wf�,o��F�M�߫��'��A�֩�tl,���1��{MGnn, y^^�`����#}�׏�`��y����l�.W�khJF48l�����\\�?.�b9o����A�;�����	8n�^�����j��)�4/��R�^��Xji���U�	H�y��>����,P(S�����><��{e��}���wv��N�6���f�5�ݮ���O!�}B�)s o�R�o���n�o��i�]��JM�
����Y����U���'�`۱��gqO�u�m%��>���5�Z�� EC`x�v���ό2䴱����:��{�h�d�ٰ,?��)`��r	����A�G��em���#�\<N��#�<?Cl=~=���4� �uDy�s�}|&����1�l�W���Z���'��/槣��[�@k���5eqV��u�b���O��բh�w�����&�:����j��+đIغ"d<M�/�c�!��P���:l2DN:��,�j�L���v��|o9)��T5C��������i�y��4Ij����v����x% �Y���sf�ݵd�Ð��Ѯ����`��Sl���{N׍���PR~'�F���C����cC�W!Hh-Q�~����x����`��鬾n,��ťF��P��<ֆ,B,��E���ڗ/��8�k��{��1W@��F�X�Z{��������4��l����[�Z9��X�~M�b^�}-��<��'�;�7�:��O�<��k}��B8��m:%e�����\��Qj���o��� 5łw4��f����4�P�}��|���]��GT��{1Le%��X��X<UNx�5���!A����/����(J��y����|�"�5�2鸆�n]���$/�s54�o�Z{��ۺ�.���G�o�Y�c�X[-�\��py��ZX��c �0�mR���o�`ܦ�ϻA5I��u��9lOj��O��v$���/ݑ0�g��1���!v.��������k�h4��p������L�(�L�]Q��CE��}M��k(�=�cwX�n��:���}W\�_I�,���R����Mm��I�v�&��@8�Ҟ:�`�&27k�>H:6�XB̈́>Q�ZE�lգ-W"��|��Պ�x��&�Q������G����vޙO�鈙��ښ�%p�%�I�p�~�}��<ex�����-���ک����	;S'���s�C2��S���@�����]�։:Y���^�;�A�<��s@oݝ�����@2�g�4���\����]��]u�kL��l�v^�A"8{P��1��R�⣰�|w�_���/ޜ;e�{�f�1E�v1{U�Yp���Ô����ddLR��{[�t�3�\�Y���)�*%�����O^ݠ���X*�F6���	R���5±2�e )�LJnM��3{�+�6O"_�xj���zs��{��Q��t�7׌���^��oq:�ͼq��W�E�~���O\ތ�ǂ�����-����6���d�PV�%� z�z3�1�b�����	�kk+��~�-w^��2a�?��wE���v�"�����(G�4c�I=i2~���d4���1K�l��Xk�m˱q���ON�xh�2O0�_C�?U���bw�k\e٠�����o����'�
r]R��dx���bA�
VO��G2����N	���� ��ss3�=r�V$Q?���w���/��W�c&!���;�eFjFB_b��P\�K4�z~P��w�^����;�	,k��M�0�m�B�0���-�e����I��4"�b����xu��֮b�~T;B�o�n��F������3^��]��ݛ'�ڿ4�ԓF�≙n�oYF�lH_��r�nrp��՟N7S�Y�!..e�Y��_��Ζ��[w;>1���%�%@!I��ve�B�9P���}ߠ���Kn�L�3�=��FԸ����=o|W����[�Ҧ2���g�_�t6�@� "B�K�����y�����{��{��M��m߈�ea`7њ$TOL ��5|����}���B�:�Z�.y�a�t�>"�ʕ��
��>>Rͥ��XS�߬r0=��И�T������[)V�j_��o$z�Q���q�����oH� '<fF���d�w4�V�CŐx�qJ_;|oV?��y�\yo�λ����@���L¿��+$��tZX�����d�CZ�u�3h���*W;Q���T<@�4�o�z�M��VU�`ef�q��
��'v�X����.r��z�A}�.W*\�c��Ј��۶�(:�Y�v����h��;�_��ɆN8)0���d/
�thyt<�O^ؔ]Ԡ�so��m(htU�J�*j�T�%��K�YQ�T��E+n�/�V�Xq�]}�f�)���� H���5~�xh�4	�ǧ�h0�ģ�8�P���Jf�T
�J�Α�Gk>gpdC�����	ŕ9����G�u̾�<-OHBB�g�v�V �pӲ����5�'�歕�E����i���-,�v�*��qm�Vc)��YF��u*�Pjݷ��&�V��(�()�%���(x���iF���Wʷ�߶Q%���N�Q�۰)V�]�9j�O�%��R�Y�=~��2��)r����"����B�72l|���s^���\<�{HZ��&TZ8 ?�H����v���6��}�#w�i� &pO��,-�ߦB\��;A܊��k/l,y��'��:Y���[2��Tq�<�7�=�e1�0k�뛲vBd/bT/�ǮV}!��O�uԏN������yp�rձ�$�=�r> ��3��ȼ���Hjw��h%t�G�vt��KLo>N^�L�����8���{�a0�L�+#Kp�;b��a��sU��Φ���7tP�����Wm���Uj�� �?O¤)Mg�9,�4��F'�u��[\���0TS�/W�O���a[�0ػ(�z��|��\�Ŵ���5�(���`��r����ژ[!z�����bp,��zI�P�J1qLM���r��u�귣�Yw�Φ��1�yO��  �.x��g���A��q2�o�u��&������B���=̷������#�+�+�S�wK�t�{�e������b=ac�	323��/� �S)��нt���{��y�1I]!8.��^Tc�<E�)��|�ꊻaz�5.vP�A��cp��L����g;.�tܶw�?�mL��v�R�����:�����{�����$v����Q䢪�;-�v��Fz�%��|��Of��.�V%�V�/���0t��P��*^��h_+*'T�8ˏ�qu��.����x1_ΨW�8�߳HA|�x\��mĜ�Ɋ����fW�.GGk/�g��8�j��{I�~@"�d߱�C���.$ҹ��q{���bZN�;�/쉼x�8�r�Z��%����YS��V�����&��<v܏����Zt���ܷ[��	�DPk$n
��D��.�� z3��Y��%���J)h��֣�K�K�ŋhy�n^�������|�c����w�2՟K�g!�f��ЧD8�;��be�����I���x�����CO�2�|��^�Ѧti^��a.A6�2�:��US���^ɖ ��S�hG����龜��O�/�~����Pb1��I��8^���z³Iwß���-�l2S��.�$�$�)����6�����n��R2��'n�;�z[_y~/�<��Ėe�=��׻h��/���yf+a�O�\�U�+L�P��T�
ʻ�?FYHkwk�m��It�g[������t�!is��R����M�<��[}�3�Y�O<�;�����X��C��7��KK����c۶��fcӐ�L�Դ��~Y� �/%���Y�-�v�]q3������z��/���^��	A�4���;v��owq=q`�aht^�n�gygɀ�qٹ����'�&�����ީb�H؋K�ÚG-�
־�1${Yi�Oe���Y�^38&Ѣ���zVń���=�{�t���fS�iT�hO~�H�e���J�aQ<�*	u�}ы��O��4���	$*�3��]��M棌�'�tj}�3ro�ɊG�ݩ�I!}�b;�֌�,�?��S.�X���B^Hg �ubZ��QC�4V����
�,P��q�i��d0�nh�����}���GU<�MB�^i6��%B5/��9�Y�����^��.����}<[����q�A:&D�m5�cJ1޾�V�6B�I� �P��;fc#ҥUOL��/����2Ƣ��ǋ��:��p}��5��SS�#������q�ˑ y���Vȿ���G���nY]L���#%~F��+�C�0�n���'�j�S$��Q��C��*6�^�}�0D�3��۫WP�6�ar/���}�f�$���%����	~L@�ג�B�Ĉ���;�;�[����w��E�"�D�ѣw!"���{�=z'��[��F/c�}��������-���Y{���>�L�z�	ŭ{6��.?��R͐f3j�(�4�\�����XtP
2������q+30p�"R���,=��R����LѮ�ZY�T��ʿV.{��8Y���_������d�n=��[�f\��ֿ�l� ��צ���Ƒ�9�ƽ2�h�NW���ȹ���n��JW�,>)<oǛ?�{m��feK<+cb�nB�_�38���m1,�Y~��Gn�a�{KⰐRF�'曞������3v�'���&�JmseS?����r��ɏU��Ķp}/&d�[JԸ#[�=5�dzWfF�=>��42(���ڨUd��9�����ӻD�M�K��ۂ$C�he�N�g�L�`U�=�ȏ���끠�ga��~�EY�E�݊���`���ۯ��t[�����d\ĉtoe��K��/=�B^n�7��� O4�O�Nh`{����B������%Ո�3��J�Q��La��Jg��o�L���|M/�}�\�G5����NNƒ�� ���t�*�|U�μ�1;&�uM���Vs�l�g����N5����1`���B�z4 <8^��\$o,.�z���wk&��z�'�_�[���P�z�R{�<����u���[n��U��ˏGl�v����I}�i�y�t^g�lp�Jz,��Ĩ�����Ϟ5��=�nsv��|���x�CJ7�Z�%$�"�ȁU5��4T�g����@��[�H��p�PH( ]�!0�E#�l���eY9�b����m���WX�ԩ� n�������7�z]�#4v����~��4Tuass�ig|VE˟Dl�_���n�����]�r\��n�����t<���BC;7pGS�4���|݈�S�N�HĂ#�#68�)�ڐWSE�E���b�J��K������c ��
��������6��d��H�9�B�Ĩ-�q��.���tI��kf"2l�te�G�A���"��i�Uj����29�V0�+C���!��&���&R�gMLLp!|H��D�68<.��z�iCd����Q��Y�h?�/o�n�9��{��$��(L ���3b�\֢7\Hf���ڦvE��e8��G<�� y�ҋ�ǻ��SX�eH�d-IA��yeͬ��2,����#WS">C�v�Uho;�}H�bUC�T	�e�h�拴��Ԛ�.փJ�U�4�o�+u�=�pk��@�^�%n�)c�5�pl�n�"(�n@�%���sj�(,�tu\)���
��[i�����������3��y�j�W�b
�P��op�8�m�"�r���v0�*����T��?�p��\���|�}��P=O���c�����D���^1+f�����}�?�v���4������ٵ��}ruРi�BE�cD���rSx�db�k%zsY[i���^��6õ��4KϠ���V��sł�ym4��D��v���H�T,��E�(�V�4�Z��ش46���s�~3F�,k*��^s< ��'�&!!��keOeUdx���eW��\�rQ�]I�?=y�?��b��o	
n/��t�fT���7^{��T�T�jN�Q'�4@��q�����`rH�1�_f�����Lv*3�- 0�឵)�q�@��֓\�1��q��ZV�M�����eVsᔑÔ��՚��X�v�DĜ�y��gdv�n?�*�I��d|�vv�~9�lXx�s@L���ͤ'9$�M�5��Hз�])U��uA�6#���Mo$q��,�;��sʇ�.�ί�ƀ��O_7��`��6����@�h�6��g���[��T#��>��x�]�vx#
���߼@w�K�Wgu��7��K�vu(*�f�_�7�o��?`�b�%m��%�C�W_��-^�gs���胏t�-u���o��rB��T��sƋ�qUʋ�}����Y�����e�O�@��H,3�՘o9�����Q����+jM���=��v¸U�V�N#�O1E�qw�w����}�	��-=<���r��n+6I���^�s���W��I���&��H�lOd�?���Y�9R)*`�艸�b�*��P�=�i��l�LN���B��I�)�YM��[�]�I�-����ڦq�Ux�e�z�|�'+%p��P������4����\��oД��lLc�Ot1(��CI�X,`�x]�.�ۺ�?��+	��4�?����TE���s勵�0d�D�[r�`�����o=tv!�Jm�Z�~�~gE*婏5��j>�|
�]yj;ln�_`8Ϙ��;����n�F"�W�t��(�-i�1��l�jBU?Ł��l��3t�}_���h�*�����R�$��ɐ�-�z��+4����|H?���mD��n-���Ǣ�%����31*���6�vb;�kb�Lۈ�-�����e�������\_Z�촗�c[��I	�����&K��@���C�3�\_�i��dҜ����:[m��uI���50�6v�( y.�h�rٵ��A����ӥG w�	��I��V�_u��|��  ���h��(ea�#�C�ɱ��)C��F�Tz��Һ����ֽ@�h����
�'~�/e*{k?ҡ2�B���S/[@=��~܏~��2)�^������4c��,Z���#M&�d�ճ��A��HNw(��c��J"�}��r�����A�FC[[�j1�`�F-g;�8����?Ɂ=�_��nZ�����҅$�F����r��d(?�Y��ډn�֩gA��ԇ�䷌�;=�J��S�'���:v���0-JSo����~���������������I9�2�cC�u��G:q�}n�Is�nO�l����5�J#�Ȅ��F|8gɇs>\�*�~>��&p]klo�"����I�Gƺ]�q=�ʃ�����vC�D���s��Ƶ� $ �S�� ����B�B'�bj32P��F)�eD�ì�g-�wv���>F7�U��G �Y-zn6�<����0��[��#{�>���Z/V�A���o�B�:�Z��鿹��R՘���:�)�m�P����5�����O��5�����^��I���a�,��VJ8ո��
�b��J,(�y�������J�V�����ż��6�)F��H߄��4x��J�$��?��o�y�(=m���f`�^w�>:���b�BwD|~ ��A]P_���, y����V9SkGA/������0�Ӽ���È�Qw�+>P澠��� �8]�U��x���T�L�����i�oX�N-����������`�.��0���k[���'��O���.=�~5��������=�md���Q�U-��y�_�ʵ�h
BJ�6�=n)D�G�Yq7		�ns�}y$�I994�x��)e" ݝ����q�����ɱ�ѭA�#���gjb�uE�M���ۺ.�dBP�#�[��S�:����h�fO9;�$�w�]&No�ѹs�:�9�?�j3�I���[Ѽ�����C������&w|���X��4�w�ݳ�i{%WIwoN����[��}n	�?
�Xl��iOt�4�>�{_���f��؜��������24��a�5���|��e2����pL���!�)9ws~�M$QJ�VO<�@���q#�d�'=��X��bΚN��Y5H�����I1F~Ό�x�K��Y��-sX�8�KD[\p�G�X?�i��NH�/��uH�ʿp5*���{k����ZZ�l2"�Q��s��$��|�g&~x^�W��5���SXID��]6��7��� ��㒹�D	>�P_�|Z�0�|��^���E�8u��X�]@k@v\�l�ȗ�:����U u�2�Xw_9ġk6N
S��`��Ñ7�wwv�l�S�k�'��3³�s�k����+g{p���qk�N�ұ|���B����U���f&��蝧�~Qق��p�&�&h�p�
ם"]�����0��!f��'��d���5����Qː!�՞���9c��'OwQ<:�:o���z����ٹ�(9� h���K�ګ/~k��%c_H��+�?�\L$��%�Ӹ�`֍-mb�"#.3��f��;��ll-�Pb���~!�>�3���È3o&\�㗸V�X�-�o���eLvr��.F � ��IO������B2�7ݡ���";��|���z��
l7��򚵂6p���}���V��?)��D< b�\��:}4ҨdN?��	�*���L�K~��h�o��	61.v�4 ��� X"Q[��n}��K�:�?��^��zR�\��D����6O^B�AM5U�)�,P��)�T�Q�劜�NJ�n�Ϡ��`i��������4/���啨��]z��a��� D
�;��IQ�P�a��%h\��Iۈ�o��� �4�n=���y9x��kva�u�M�� �Q�އw����+�r��X����e�l�:�`���~�a��AV���	H6�he.@���>stw�^���o#FE��K+a����;�&�_HW�[�ܪ*�����2"�W�P&	LT2/�/kg�N����L������H�������D��T4�v,)��B��Ue<�+=�����޹��%��^HMd`d��S�0�?�ʂ6��h��y��T��ʝtk������uQ�c�v`$�-ٟ�O`�fP	)���(���Y�|)������!"�dp�F5>���]� �m�K��߄'ʰ�v�����a5P����`O5����/ҷs�S5��M�r;d�+6H�(���v�0Qx�]3v*]�Ov��SUX���+�En���c�%B���}Vh�rb��ڭ<�' �T���⁛�ҵw�AF�M=g߳7�.��y���D\�}*A�##������/��O�V����-��z�E�E)9��m1�+�1��`�v�F7������+�Mcc.�,N�rDY��
:��5Ʀ���8�x�,�7�̒�9�|���,�OǍ�EEE뼳�+�m9( ���-<��Tm�`6�~�:sN	�Q��ڵe���r�Ly��pm�c)�E>�lr?'�=�o4_��H��a�ʜ��l#�)�*d �7ӵ�Y)e�Z�v_p�i:�rH"�.kH��~���]1WX�|g��NI�	�̢w��S�Wr���oc'e)�x�[�*;B�6�,�y���DH��mIm���#�{������T�k���T�>'��Y�4�{��15PۤE��ҷ�~_�������Q�+Sg��fS�L!U-OC����1�D2(曢�L��7�����iL��u?<��i��6�R���:�hJ�Jګ�0^���AH�6�
�C�`JCkHx^t�Z��OM�b���Ѭm�C}�/ck5F[���3�t+�<��}
[�5��Wn���_��ZO0��H$��W�l]爹p������b�񢹟msmV�n,ck}�,c��ײ�<���Q"�O���ta�"�c|�/��(�D���Ϟ"z��x9�[�o�!�iu�wXX-��Ӑ�����e�k�oCεr���{������dܳ�?���B��P�sT'�:i[zQ0�տs�\��*e��9J�A֦N���GY9�S/R�>h���w��qx�j�M�dC�
�n�������qe�$|S�Y�5���_�So��	6}��{5��䰖�br�ӝZ��?� �_FD�3g׾�]4瘜�Cש,mE]DR&��8%-��j�܊�m�����sp��CW,
5�J�Z�)'�ͭ~tP�/�k��;Bޝ�����-�)+�z��T�����-Z5����#/M��K�JWf`������g�z��K���_췮K~���4�i�9ih�������# ������8���ZK��#}���}��CB�>O�v!(|�(e
�@Шe}[��)�y}ޤϠ�"�?�d�\��Ǭ�)�'�p[_z�@�X����;5|+��ʜU�W��y�M���'�e0��{�>�j�(�?v���&����֪E�R�R}���T@�t��R�B����e2.%J��A�2��,�XJ��,�Z�.�o4MR2�������R�!���G��]��M�Wj=�Jl���6�]$�7}�'H�4bԖXR�[a�X{Nh:	L���AW�4G�4x{xE/fS���Z�ڣ��ipØwPYڮ�*~���l�M��c$~�D�XO�;ZKÄ�9&���z�J��q�	_��.܉h���0���а�j��-"A�!vqܹ�q�P}��|�+�<�s#�_M�}
>�9nɉ�2�^4�Q���,g�G�����H�ո����.x~8�o?�k��4�JE�
�R�2>'���u������0?��$| ��R�_2a�BU0������.vZ/�u}Єe8@�O���O;k��G��?=�}�w��	�h3ř�w>�	h1�KC���4�7��-��q|t1�!���w��[u�����ཟ�%������2f��(�{��b'X��N�˵�-�x�b+c̸��H��,�\t�6P/>.��W�kf�>�3���|\s$��g�g:(�0v$I���@Ov��5I%TfՆ�Oz���^���xws@�'�|���e�W�B���P���X�� ��$���]s��?SUIJ�.1��%���X�,Z�\���x �y(��F�`�WVz�|W�Ÿy�7+�/9�n��j)i>��t�݄h�w�TZ~Ͻ��Ѧ�w���?�Ȍ��ޚ�i�&�-Ɯ}�'�ݠ}Y~+��z%k����_��B+�I�R�+	|ph	�9�䋌C�l�@�N^�\>�X�p8�o�z��D@�ƝT��T�������0�`!u4rβekC�6�P��w�	�L���ս͸���Ƞ%��y-�OB� ��`�ѡ�-��n��2��v�V�克��xc��ϔ��=S�?\��B���61��V�zvQ�q¹x��oL����tG�I��-^r�����F��H�e�G+N��Vw!I�YzϷ��76���S���� �(DQ<_�圁��Ӌ�bf�P[�D:Y� Qo;;���FcR>�һ�
�njA��f�fK3S���84t�>s+���$�<�������w*�n8/�~��b� _���K`�*T��=+D��$�tm�HC���x�\�;��F���~ya�B�,����-v��Y/�r��z	��{�9��׈E���q�Df�=���B�Ɛ ;Na��B0����kA;	\��?Xm�]>�� �2<�]��ą���c�LI���H��ľ^�����r!a��W�.��$k�8��AiY����x��d�.�TDeV�!�����율�o��S!;�� �_�|ꆚeJ
�+�ѱZ9l�_x�b�����S}'��<�����B�H|��u�G9�����;��X�?]�*���jy�'Z#��s��F|MzS���y,�.�j�Ԩ�r��C>'��Yb��0���ۏ�闏�/�����~�
Z�J���+|���������	!f�J��q��=[�.��#���!�����A�|�> �8��C��f2�gZU��$W���-�7U�.[S��з�k�N��t�����" lkT=����cM����~� ���AHh_���F��,��ZzN����c���ٚ�:���_�ݖC���xX/QG���������n��EE�����F�ꑿ�:�'��I��+:��.�|��=�����/��Z �h|���ى,���|�Z��7��7Ue�}��4�<��N��}�z��_���E���9d8� ݍХM2x���#&W,������Ai�?>�Q�ώ�=��&6���
�V�._��_b4v���d��k��5��S�"�޹{�d߀ف��d�
`��)Fj�i~zr4Ƹ
�1�ݷSƙ(������O�Bd�s��nB�c��"�X�O�lTE{���+i�*IV�\�����_�7�ͧ!�� ϸh�/n�X���͗G��u���Z:!2{��Ih�@���A��������D�o�vç��� �6.c��?q�'�Xtp>����Zε�(��M�X��J��V�QZ����r��&%X�)ɕĸ3f��~�/����������d�N��wך �y�+;*vb�r�2�M	�|v��Q�|����R�^p?Y-�P�6F��JY���!~\Ր6�>HÕ`��l���4uJ���Fv�'�r'5���nz�a�O�ō��R[��������W�L�3�ZV#8R�$�ָh�j�T���:�q���{Թ�y�r���K���_3���礦vLh��y��Vt��.SJ�� �4��"�DЅ��a?���2LJVS��W'V�p|�z~oA/4A�S$J)��h��.0V�Yh䊟�Wq�dO�F;��8W:�a��=/�`���\s秢,�fW�v�	�e�{��@19�ZE�Jc���Q�i<xV���띶wvQl����/�^����\Hy�@^��V�Q���j߼W��㧳�M���V�oSh��T�/#\ͼ˘Z�E����c\}�׈h�����ݻ��UN��0��Y��� ��Xl疷q�X��o��;�	��s� +RtǠő;�D�z�(�hs��b$&i���XY$����T��}��ئ6��O�Μg0M�5�}$��N.���0��ߘ!�j�)G�������������j�ڶ�LeMW�E�ܾ��鍾TP��f+��;I����E�>�Є���-�E�a�������W<��gs:t�-�%r@[4g����' ��ʙQ�qk�'k��Wj��������b�m"Z�j�b������f�p_���{.�	]5�v$ǣZuv u�)�-�*~�����ܚ韜v�'W�M�w�4_���d#Vl ���B-d�-��6A�}���n�������ߢ�)㼖�Q�k��}�^WEQ���h��c� '���Á�6�j�����~Z�+rN�Y�W�Qywv��-��w�)� �֗^7��3j�C����52 �^!5�
qG�	����������{M�3�²�7S�K�$E,U�Γ��{�0EHn������N,�W���c>�~�my�Uل��7UvZT1��у����jRy�9� � ����0��ΦCZ+X��B�\.�+/�k�E\�$/;��Sq�_A��O�h����f�tX�bmYo,�Cx�qgj��+f�</��p�ĘZȧ3����h#���Yw���gZ<�q�����)���Os*�g�)������֜���5�ף�P☰R-'�h��7�d���s#�؊z���)�u��1`���k7#w����g}��K�f�Q�'M�3c�b+MՅ�H���.�R��o��3�����0��V~�7aK0#�P!��Jd6�$cPj�ġ�P"ɩz����?���{�+�E0�z���a{�-�!�pI��Q<�%�?�m��U��+("�+�����|6��"�����:�����U�9\�6��ߦ��b=l�t�a�ә����8E��\1��#�$0vp>m/��~[{m�I�d���g,ݝ�}���p���ݭ��U~����vۯ��H)��;ۦ��[��F�+�k���:v��N��2-Rƛ�����+�j8�ό����Zdה�G���>��0�Z�'�ɝup��V��{�$�B�?�ep~rx�,cb1jюr��W!#{��=�jd��xM�,{B?~��D�tFW���g���co~���m�vmp_���Ђ�u|�o{�^	_���4 ��m���l'�2..�Z�U���W<{������y�Y�-c�oa�Y���q1�j]z�#��.��ƙνJ(�͟,!Ͼ�[��>�:SDW�h&���<�^���X����/����r�̡0>�������Dم�ڃ�=[ �<k�?$wS߾�Ly<�\�t_�>�#�}����gC�4���ю�,B-l���� ���MG���)�D��9��?�-S/X<��n��& �S|ۺ��6�����
433����N��<���vq*&eH�B������G)��!I�]Q�er�ڨ&J^�M���3�7�ewL�ٚ��t�1��w&1��-�$��{
�5ބ�ym��f��	���S.s� �yY>�xOu-��=+쇳��]�Ęï�tE=X��/i�#���U]�gJ���g��{�~�k]X{�Q��sYa�iJ��^�&�B:蚦g��k��!�F[X���K��q�<�aܪ�A�^f�g�5���G�������i�6��"U%`��'��u��蹵�+I�I�s
�����@�y�F5��-�T�t������k�rO@?���qyM�U���e���F��P8�S,�h�52��MzAc�5]����(˻@����BӅ�dh���D��6���y#r����)������(�*�>�vs�!bV��w����Bu�p����`Z��"�kf�9dx�D�Q$y$u*7��f΋����E�k+(�x�8�t�h�*��V��h�?Y���c�;����$yeV��B��j�i���Y�^�;�h�j�o�n�V�liޮ1q})��
ʇ�zm&�]����Ō{�y��+q��N�-�=Fz�)/�q����k���ȍ��>�q-#UK$}����|�fNkk?�֜匼=�O<�vU��۾RbwP�Wl<�HE�PG��ߏ�S~Q�#cףtLf�1���F-�\�7��K
�sU*�F�{j=Ł�ؔ��.1������G��$?&����'�b�o'�Z���z��6�����[Ѩ��~�n�@4�ܱf&��Ѧ`��?�0��wNEoyq�әU���v�[<\O!��q�7�U�(���p��_�#9t\�#�VR��r0��⨻����З�)������s���S��������uQo�������Ep�6�wm�2�v1�R� Tf<�q�k����9l񳫆�RJx6E8��s�ra���b�\H9L�y�cQT�u~��N�݉������*�9p�
l�I!�K�-S��q�hق��et�4l�Ҏ�����>��4�Mcщ�~�����R�G�ti��ݼ����u�V���_ż���A3�oe���Y%�5�5���i;�\�j�7E�G�";�����Rߝ�����v���\��֓?np��;��dv��k��B/߂�&_Yu��y.Gql;���߶�Qʳ�/�g�OEhS\���F�N��\M�1�e~;���2�g�k��#JJ_G-Cjʱ�4�/��~.�;J"�g1�hz��$c��J}L�:�o�a�b��NTYy�qL5*_#��� �c���Q9Yq'y�ǢhV�,�ϰ��S�� ��g�oy�(#3��w�9���v���E�s����=ǉ_h��N4E��D������yF>�����.��$Ei�Ntv��E �K���{4~� 0�T2�k��x�C��[�ĩM�0N�ߡn�3���3�;��e ���� >å�#�_}��dr�ᮖ��He�FEDR�)]�����޺�)��-�	B�+[��hֲ�̿ �Z��T,�����e�b�.�0�-)ꥃ�fk�ʜ6t8�9���*33��������`�H/YmW�Q�y_���n!�KϚ�~SJێPR}!k�O��MU��s�+r4��待��5���:��i���͡���t��^��W���\|y�u<�'4-��Xu��gF�ݲ�?����?XZ�C�`	�kC@.�w�4��s�%%��������8J���߬�žMp��hԶ/���ۆPh�;��V�I	pb��Y"l��k����|ƨ�<�pe���5��cDX~^�����!'��3����l��:@"���rؑ�|
�D˟jg��5��oXI�ڏ�38=}�W���%6�%�n��d޴7΅���ϞL�j��������,�mV��,N�lj�a�g�g�b@���3�M��Lj�K��Tm�>�\PO�0Y<I��[g�b5�pC��l����W��γ�Y�EQ�����o���/���9�2������������	
�Ʀ�
d����M�������:����5����$��� �/�>R�T�ʬ΃s������`K՞����a�0����}_�N�i��#��q��J��j&���`!����?`nF��l��
��N�4n)A*�@�,#X$7r����y-��;ڼm��Ͽ�Qn�|�4C�D��q��>C�R������Y1%���{=��NQ��=�&�G��Hs/e�oCD�"���t��dY�@�����o���q�L��!ô�&)�d��$��Z��O>J;���j�%?�V�2���WK�G}��39U�$b���7��J�K;��3�*J���0���d���0����ѧ���ҔUɣ�|3��Qӧk�=�J1�a����b��kM�>Nۣt�35@�*��a%4���R�?�j��o�b��қL#ۓ��"��\��Xr����
���=n>O��?Ua�[~z��������A���?&�����"v�5.Q���iGgaL��9B�֣��������������ڙ� 9��ICߢǜ�A��u�;�{9�[A�����%��_S��l�Q`�~��<��~@ŐP^������ރ�|�>�-���0]j�V":J�>�1�D=�����zcWi��J*ɢ�?ev8��x�Ȟ� �܋��~7��CţTv]w��ǼBufrR�3݊$�:�{ު���%\V�Hx��>�O��`�W� �Fy��3�t�+v�r���^1�V�X�=�������K3��ip����9BNhJWo��<�
��̇)����;�\��~�I��ʇ����)�,�S�F<oob���T?{~�B.#�r���U�d�͎	G��y.궸F��IR��C���e}�nt�T�y�b^�̪�I���x�H!�u����+�U�t��h>I��5Z������U3}kQ�"�r�*@VL������4x�-��v�ٳkK�*Z��F'5��g�~ɟ�UZ}�B�%��lKx��^ϒ'T�k����%nDK-��:��X�4NK�#5{%2���J����D��-3/�{N
�g茒�s(��Z^qMv�;����Wq�7f���r�V�27��ˤ�_�뙮����<��Ԫ���<BR�H>�w��VP�����L���{�.���e���f�'������a;-��+�}���|s�
�AVwg,�4�
���b���bn�*�m�)�~AՅ�2)�\��1�61�޺���z0CE)'����X<��>���`/��i=.ģ��tSn����8w�t���Dx�'���%��*�շ�n�i����2��8�Ü���V��D�
��n]1��V"6��i�om�!/�[��.�JI�)yn��v�2��iQX�?��mV��L��G��J���p3iS�c����xw2H姄D6��Y��]#��KVB�Ҡ^LSxrày�uD��.�L�������ݫ�ے��MLx�!�k%��%Էy�)�ft��bFxChVƪHG�K��dr����8�Q�a�K�J+��2 ��_sq���;d��gޙ���r<W����eO���pEI��>�b�آp�ĉ�mW���(K^���Yݴbҵ+1~pL�c^�{ʫZ>c�'��?n������v�=��4�DHJ�֐�a��Ji+��nZK�_�g��������BAm��_����~7�F���)m�>M��+0GNӨ$�����VN�.4/������oWV������kCj=#����E�.�!T-N�{�Z��E�Z':��������.���ǅ���%gh�%H����,*��D��8�}�����K���� ��S|�o@�B�ʔ�c���i&0e
й;�1~��;.�&�*��^��}s$�;	�P3wr)+�0]�g��IZ4�s�Tkxz���ϭN��������c�[����p�8w߷�
Y���]h���4����I�J���hգNك��i�I�������G"�6��2�ߵ��=��7��e�����W�B��0�9��7;�x!J���QH3a�K�	�NR���G�P������o/��D��$�)��=�L/,Z1ʕ��(Kۈ��(C�7����HD�=«P��85���9���VU)�j̮��&1� ��j����FCo[~
n0>s��������v�dq�ܻu�Q�N�AP��7��
������ybب!��[�8�&*h�d7�5�ػ5�!�gL��z)�ϸfx�#�]��5lԪ>���W�[y��M^�-/�������\\��y������-V�v����>D����,'^Y�omܦ��UzVa�~$R�Plf�DA�$p��#��k@��}3!|���#�>n@���S�Z$'ٷV��(z���TJ��@����]�	r�w�gM�*#�`2���~���B)�Ce��5V��nZҢouY/��t
�gn��>���Q����������G�Pأ)���vz:\�M-�Vs�u�;����N�j��a�ۈڅ����A�V_�M����V�cة�hZ �o9��݂�H��RXg��$(�41���rz�Q��C� ��~��G�KK7�2_��9��sLN��7)�y�H��c��7��wC������yao�خ���$k��y(Ę�Zߏ�M��g ³�#7�=c���o	��5#�͎��a���5�6L7�hk�k��WX~�����Y�3qgm2>�0�ؙ���!y����u�83֌68��o��{���6,D�L��r$��|�< U�|���
Q�!�>�7�G:����į�>;��,y֤ăX��r���j��4��ΰ�����TV0�~#��^�+���k=]�hoԋG���f@&���J���eԔ�h�=����~5��O.��ᐼe��1^��y#m�H�{���N��Ѐ	�P�����	�U���B����\�3L��Z)>,���眏W��%�Q^+��X��������k�V���̄����$NX�q-��_�g�S�&-=*1è����%Q�ä��z{x�x1r��Q�w�l�����芡ꮌZ�y04ؗ���;��^9{�k������[����&�H`[T"9]n���\�K�o�,Q;�t��M�iY��¨�n/&��������"E�z�����;c몿 ��.H.N0��C;lM6;���Eo"�e�����|ޓ�l����o9��
�����, ;R�H�vl�[����2��;�9��g�Տ�������3�X��CCN��Q��)����5W�f�>��ǩ�	�Fi�$YG_��C��s��BQ�,�v>�w��)g�_s*U ���aΝ��:�/�S/��^^�NY�;4���g�,;���
�m.NR�K[O#�� ���>KO�Y�];�Ӟ0�l&ȹ�g
���Y:P��<��^E<�H9i5���4����������~�E���[wQ2��7љg���n�υ��͸L`M��7�-��?���&8+���o/�0�d3r��3��̓K�_���'�y�ˠ���x��v���rl��s��O����ވb%�!�B���w�CPB˲��/U�q���܈.�dTS��RWbՠ��._�u��9w�͵d=�J�i>��p=��4��4�<Oȹ5�G���$`�<�$zjl�gQ�����q{9���ʉ��M�3���!VG�t%�Jԋ�K�%�7"�o�ká�'��֯�*Q�~`��[���[�p�H
bU�_?���\+Iu�Y!����4}굶�<� r����z�8吤爋U ��3���ڍ9O�#�6�>F���A� �=1�`�^�cxV�0�ү�մ�QD��ȑ��P� ɢ��.��o��vL��0ߓC7�J?5�BC:��x��>$��c�|��>��Cβ���?c�U5!p�N���B��ܜ�[$�W�W��?��ۢy��I��;r��̆8��k�7�uD������}1Z���"��9�1�O��sMa�� ��zz�&\4=%�A�H��1O����������^�z��߄[�k�2ȿT�C$G�N����֋�J1W%�qՇ���*�FvP�Q#'�r��
~Y~,R�#��;�C֍Σ�sR���H%����=��`)h�Qf�,N?�Z��_'{�/2�냝��̂o��f�O����q��Ak��"}���/6���X���R�}�"�of�Gz�����S6�I@#�\��K˽~�I헕6b�=�/G��JpTX��וk_WnI<�,�+�o��$�sYQK=����,�F%���u�x\��s���� ;kB����ny�em���^\ y�!�Z���U+c��z=��P����~��Kh$����֒Әf��%L��?Ը8�i�6�o���w#�	c|8�Xw)�'��7yE���H���&��w�%)��,�N���2��!\w��P�]Kv�����%���͍%NK��l#vQV�Q-�N��0����p�\�T~���z뇦��{X�iF���[�n�Na�]#JH��tw��1P����F7_�����/�p�s�s���3�"�� N�{.���nP��G D|��I��4MX��k��~�F�vo�<ϧ$y_���Ud�ԦX��V�М���4���5�>eE��Q�u=�H�f�Ņy��k@��f���I��T)Ѱ��{��X���ё�M|u�Y���M��	ay�è�/�˙#���=[���X�.�h�K���j�U"V_��.?��;jE|�X�,�0c�!�Ph̑��t�Z����#�B����<��Ӓ��>x!@�ae ��ý��%6�È����t�\��4'�7c��d�}���_����q�+A�jUU-�Vs��8G��T&���7�(j������h�|������χɹ��Zvx��ɺ�O�t��Z���� \tZ؂7�D��ᲁ/�-�����p��I겳�lJ�u{(�n}?�z��K��=��'�DbUٌ�XE
��&���p;I���P	�;$���>�R���޻��V��Ǹ��Ʀ.9
i+֌�����l&
��C���-a�u�xD�Ԣp��J9�u8�J�p���˴��W���ᷧ-Nˑ��ǣ[V=e������&`� �IkT9�yBC��*s'*j�ĝ�^�-,��*�P�I]qss�:�gu^��s���G����G���.�(ށʴ�����;�*tm�p�#o��w��P�N�ԋ�bG�)� S.e���MI;���CT�oqor���uj�15&�ɚ�]'��a𴆜&�`����`J���#4���v����������a�j���Id$W���(��"	/��½hg��>���������=zdS2��̨D��O��BBy�_|��FZ�&O�T-�x�E���=�����Df��L�&e6qStf}]��"�2�ʎ[��%�j�v\#�[�/.4�G	���TGG	{���V���FP���ӭ��1>+h�)d�e�۽���S��pt�=�`�k��&����*y��7��E��r�}����ӥX̦⅟����F���˦Di���&){ևlO�hO�QY��v��i�HP��ti}GA���	�HnM�T%� 1�9oE��0U��u%WjjZS���O���c��]M�ȳx�ߌ�����ᴌh�	c���#�v�}��/�?R��.�(I7��RQ�����2�5��*a�t�P�lL���ш�lQ��i~.�Y�c�N�l�j�U*k�ekwD����.�sc���O�:���" �[�g+�XU��沞}[���B+�י��F�p�����g���Q�;�D.��&��~i�1�����~�%����i�z�"�C(�]�[/�[>q�������	�my���)�G�<C+�:QݞYgI���y�}r� �z��3齥J���0�x��=2�u��x�wH5�8��F�><P2���w�����Q���a���!�?6�.i���b�5Ϊ�+��#�nM����`T�4�e-ί�����E^_����II8%C�E/�no�
Wj|�E#y{9{�J;�C����]��/��ݹ�21>@��tV�����8{W�/\�:÷e_��c��
? \yz��)"Q���ۣZ^I�1�7A�TO�=:��\�2��E�^���O����6�Z#',?�=4�L<�C��w?h�m�/���+���?3�f�Z�D����?/y��`;(Ҷ��w�\p��Ti �w9=M˶J��Ѽ
hȴ��U��S��L�)�'ҁ5MQ۸ah�^���Aoې��I���\dY����o�s� �W�5�!3��#�U�E�5���π��cEɜy��1_�'�m�ތ���P�����YU(`%��/�$vn�d�>���{�����[B���m��Up���������]�LϽ��/�Z�����:������B9g
�������aa9�l�U�a�+����v�)�ܲf�{�*�@����Kbާ��Y�S�4���V�EY�[�
��$^�'������36GP����n/q�7+����<J�R3�?Jҭ����v��/�}z�a�k��GV���1��|��n����Rv�^���D���a��7��lRҰ�6��z�z7�a&��q!��,��qd�N��k�2�j�//��d���*��$�������j���9���cY�z�5 �M0�f�cRE�����s�2~���t�Ƃ�X�`- Q���?��w�z�.;?��v~��v0�*6�!Z,/{&c���E,�&�c�*���F
wClT̿�²�x�n(*�,�a���F�(XC��l�nK~}�+P+�筨S�Kb^k����	h�#@�W���Ϗ��Qŵ���Y�r���SN6&�/I�S��J����h��/qT^���_��BH�����̋?�	�;k)����'zߧn��jN�x7��6�����3�]�M�v��V�X��Xݤj�l}nt�"�PN}�u4k��ELj��Cg�	�����j�#���/>(K�v��ɥOX�;<����u�j���N�cƦݪc+Y#��Y>5ya��>.隣;!���#�j̦E��H�/���v��&S
i/�����CG��<�K��L^� l�l䣞�lb&�͍狳^�~ֳ��/�̬�
\�Ȟs.:]O��G�Vn�(��ݤg��P���;��N���pj9�-ь2>�h���[׷���07=n8��@ƭ'�)Q�]D��������XOM�S�X>�q�L�M�:ڞ
��JS%����Ex����^���!���{.,���ф:ٟm��X�ퟍ�Vͺ$��-ϥ ��<s���mD�T���T r:d�_�U�Ԫ�T���+7C9d<>U
bCĞ����(���\�R��h*|z"g_��d����O���,��^O_�g�d�<1�bE�S7xL4q�U�;�׵_n�M�-^�m�lUH.L[�Oư�����O^�'P�'(���Q5��%��ίA���'ޕU���yb�s��3�Y��F~,�֓V�ew�P���n�ef��s#�>�m��m�~��tƫ��L�--6�K>nj߯��Q�܁�p�h�z{��O	B·�,q����#�?��73�+&s�n咓�]���i#F�܁dR6��t�\{��Hb>���viw���a��J�^�i��A���?-����;�/�Q(�0xs.���Z�ME��j�Ir�s ��d�Qv����~d"O�CYce/9�f(�GH���d�S�C���V�>>8^��[��n�'�b�ύl�Nz��)�n��=4�K�h�	l�~k�
�-��&�/j`�B1V��`�hn�IH��Ȯ�TvPw �
y�T�M������'Y���jw������ɷ��O�<�����]�-��r�v�9����rJB4'a�`M�����p����k�Y/�M��S�|�[=<��Fp�8�ɪ���	5�A��f��

ݢ�N�[�S�,�/V��~&�a��H$Q4�P)�7�H��4[wǬƤR�Rߵ�w�ິ�s�����xi};��VN^���K��.�eJ����~�`hl�����>�烵6��ù{����i�~�4&eX��Nl�ǂ����m��'���Z��磢a]T�ĝ�����Lə ���6��!�`h}�r����7�?JުG�Co�<���������/����J��p2�#�t}m��_0"?�-M!�;_hz~gˣ'z�Lj������E6����&�,��F9 =�*��O_��c��l~�K�N�A�J�6�1�-�V���78T�%/�ڍ4+A~��Ga�t��s�O���aFYY�z��憘ם��E:`�k�K��>:�[Ll�
#l������������i�C��{�sk����c����)��TF���0\������C�^�#�loRɛ� �xy3Yg�����ES�uÒ���^���-գ�WG��{�^���τ-`��%������f��L�Q����
���8�yK���2Lm�e��`�朾'Q�1�ֺ)�ɇ��{����95B)5�͕����;����iw�Q��Y����� `�B8��[?���Ft'�w��s��K{����[\ҕ}��D>��!�"�����S�i�}Sx�M����e�3��9�
�Ҿ��<�=�Q�;0�<Vߡ� ܚ���sa�6���m=H����n%ڄ?��a7��BS�(�
� �7MS�b��;Ӻ�i��d6��>7��̪&	9��O)}���8�zE+%},P-��\:�W,�P"Z �:�#�'M���t.�Gf�)�9�Sy� )ׇMK4c�6�����q﷟1�Y?.��lP�|"�m�\P��d��y����m�Szf{P�U���L�4����C~KF��3�(և���zH�u#0�\�{�7�v���3������2UW�)�A	��?��)V�\^������T -����f~�'���Z?5���l�|:�x�9��r��}$8f[�����G G|g��xW�BfJͯa'�޲Pd�m,+�אꖳ���u� �瘬k�W�� ���{�YF���[���!g��6�ȋҀ��]o��ω��|��:�wx������v���d�~.�O#2Yt����;�	����TU�}���r9��&�1�h�z*��M�y�n��(6k�Ղ�L��"er�iM�?8����{�S�lT��r����g?n�(���*�i�䗅%T}���e=���~.eS#[?RB�w�!�L��*G��Ӏ�S7}��d���"���e̽ ��s�)X��u΄�u��r+3�Eji-~ދr�Z ��^Bb�A�}^����B��)2�D����Y�^S**�ܒ�X���4������yT������8�Ph���+j���X;���_���L>��oc�qW������Kr�+�c_J��"5[o�j�db��7b�q��ug�6m��x�n@p

�Rv�a��ס;&�<�:n������~�xN�I	?)$�I�8޸�N�:)�'����E�úz�|m�uI�),G�ܗ�J�i�=��`�,��V��6z-;Iv��ANj�Fh�(���J��@�y(B�?f�h���p	�H��&�
P,�N>�_�ݏ��h�k��u�-=����9�7�Ϝ��5�^�x��Z��Pˇ?v/!��9�C'�s���o�d���"���y*��v&� ���i�^/V}����^��\P�k<��j�"~tC}�7&�v0�RQ2���J��t�Ni�x��K�7��[	�����ד=��8C���:�}���vKҪ� ӯG'x�Gk���# ��o��1�̸��TE.�>�:NYo�3>WN��'@�����G4���d��:��}.�>d����
������� "����1��2
���k*g�li��_C�:�� ��`��5"��c�<�%�A'���k���DI��jҥ�؇D���%�c�v��t.�c��-J�N)�e�i"�*6G\�T)�y���Yj��ѡ�HQ5�{�CϝIm-�l�sQvι��`k�Pk�P�]�b�ޡ}c���������(����)-d�$xj�����u�W��8/��&���/�ҜC��g�:�F�n�~�뎣�Ѷ������H2I����!�6��� ���`C#*0~*gq>��0ʨ�?�hg�m<N�x[��<~�eOOE�k�����?sOfϷ�K�H���E�SJbe^��m����d/�`U!���6�{ gZM���~�0��Ȉ�js����=�����'r\�i$�M����Mst+��b��"�!�WR���5l�ٻ`���3]E���PR�#�����:nD֩�O�MQ�HL]�1E���,Lk:�m{��N{Zm;�7#[7�����S*��>RDǦaeZ�}��vRrl��Sb�'7�Ah �Б�u ��%��4�ca��kD�i����6̖��g������*�`.���v6�i��غ���!5���W�<L��̏�{���s7N�&ӯ���wA5�d�`QTW��.���
����4���M�o-)��3&N~bm�{�&:��x%�'q�Bwq���);ƫh����_(M�a������Y�ȧ�3��_�?�����ԵFI��{�W���#�2]ƹ�����e֎��i���*&�-�ءFʸ�(�a꣄b�͠�_���"��[^ i��}uwƴ�鬻�'����eRo�|�O�o7tq�6�$����Ø"�j�cL�T�Ŏ�T�_��;mؙ�WA�����-!� �����N�����ǛO��5ǜ7ַ�+?����#����W��g��D�^<����uzV1�
��؍E�F>��:�&bRĖ��A���^ܟ����}/�n�@R����[��X���U�IQv�jX�I!��~���Z-��Laۚ9֗|O�෼?�E+�NM�>xpA�3�:������{ϨV��c��;�	n���-��9 V�.���wD�Vn\�.�P[I`~����ڼ\��L�j-LE�P��`z��c=;����W���X�������&���q��v��ֈ�5�jS�(c�`+�)�{�䒺�����c�����[����┝��-�͢wr ���Jȩ�4��	��. �COj�Q��P�dL��UuP��DW!R"^��8\�lŨo�Mϥ9�$����_ITCg2)�����9�ʴ��K�S�Lj�"�Oo�9�0�o�G�8�tw���B�9���y�^!?c-��b�s���"	;��l8YыF��ĢLn �a)��O�:�s!�t��!|�p��mr|�Rx&n��2��R��(	�z�<&H0~m��b$�$u��x��j�����'%�B��'{>n�������R5t^o���I	؁���{�QK��n�ϬVz{�9V*	iL����c��G!����e���t��᧍D�1/�����P3�k��k��ws���O#�4�<^���(�A��.�a�\��g���:�m��"�
9�Yh-]�=��0���pԦ�烨�6[���5���x :6s����k��o]�F��H n�6y����z&���-[`0qe��+y�S�3sO6R���������)R��H�<��-��yk��sGp��٠�֋쵘ssy�O�ή���d��^DƢ'u���ig���-�շ���Nj��уtn|o�e׿~F�j*t}1Wi/��؈a㛴��t��!�a3��>ݗ��@Xu5�*|���m/Fps���!��ٗ����E�Vf"ݯ��dgI1�6����+<Z6��Ao�̵��6oN��r��IFw���e&����t�T����W�KN���^�Ī�lX�RFDY�'�u`�lq��ܐg�*�Ų��������o��0���}M���'��l��ct%<�����a�e�uȘc]Ĺ�m�R�*u^��7�j&_�ꕎ.��5RU7+��`�<�ײ�D8��L2~P|���tw�,w����r�5Qҙ�8�pq��½|d��{[}��z���zAR�5�xTWr�R�ۉ�6��+.�f����{(���,�,6>:V����v��ԝ}k�Af���v�U�t���9'iΒ�>��ue�tN\xJ
e��`���6�ng&��s��w�CJ<Y��rZ���3�\�YZIx��A1ˉ�n�qO��R�m�_k�p��)�&�{p�������Ւ�.�|�����q9��V�ttlVx��Ma�����R;;���R�����l�;4�㎣�	�'�b�t��NSn�=�@��`i�^�7�0No�
mD�%֍ ~�x�L&�g�}�I=��{��(�� ��L�CXPL!���iw �;5W�b'������B?���N������Q�j	𖱵T��I�6��{œk�Np��/ׯ:1i�40�Ϥx�%$�x,�E��g��&��1Yy�'�Ӫ�O�g��7B^7B�Ŧ]���7=�D�:�5��w�f=<E�Pĕ�k��Dٷ��$�5E��\y����[e�65ktW@ŀ��#B�w"Ap�O�����n{~wی܅ŗh��[���D�{�Zwb���Ix_y�cpWJ2�G�"���Y��|#$�'o����;�L�\�!�<��Iൖ����w����Xs�-i���2����庫����Fƴ!���˚+�.O2�ڼ3�o�����E��P�]k$T����*����n�
�G<z�ώ��ٝ!�cWR��즧hfZ���&���6���[�Z�
�*����.��%o���ihK�b�����'?�����v(��ڳ|�uf�Gq�F]�ϝ@7�{m�����vL����<(���H�i��gJ�0f1�3�l62�X)=t�Ƙ�e��g-햡���B!�v�@?'���-�������H�>���w���V�[�[��Ŭ�J6^b.t��M�X�B;��Vuڜ�,��<;��1�c�+˯�b�%j��kC~�Tx��0D޹;�|�:%����d�\�0uP^L�MV�.�8=���l������5�.:[^y㠻J'=�aջ�y����rRŌ��SI�ւP�������fzA"3e_�'k̈5Om��]�j�h/�V��)P\Ȅe�:�/������ᙔ��hG`�1ﭸcۑAu~R|��90Nt��p1w��y�n�5�R]�mZj�z�����P�1��F�\�Gab��/���Z.��Yf��� I��
�{X���n޴(�I��[|A��>v�9��1v��
ˢ�mA����첤�M��)�2�2nχ7\7��]�����P%�fI�-���t>��м����@�CE�"~t�r�0��,Y{��v�d�yN^�6��f��V5mG�z�&�Q�'E�����v�Ā�]ҋ�%�����m_��rj|<�7W:d��>;F�}���9����1-*�[L�O�*"��a�����s�Us����JVz�Y�d���H��&��m��Ơ����k �m X���:������:K�In+�߬�>9���I@�{p�3s>_�_i��"4:RoW�VfV�L��h�4���7�)X%}��W�c�����-��3��i�kG��]E秧?DFL�����g��獐� �U����X�L�.�jp'/�
)s��;� 8|�Ѹ8
�J���2槹%bcnL�
p���U5V6�kra�}�W����/d���i����]�����%a[B���W՟��ߓZN#�4-4�!�Y�~����G�c�f�,x� ?
��F`��[�gqb���K�O�vD)��-��yS��f�^U:��ڽ��4���K+��݁om18��XӒ�"�:��.fЌ\bׄ\⇸�W��n�	h5�3Z֞�������b2�Qg��E����"b@)9Q{���f�C7���ּ��KiI&�3
�����Iu��u͊�%���<�M|t�Ա��� ��H.`|,�����b������e�˻�2��olB�����+b7�<���YĖ�[�	j��z6֜C����U=E5`���|�mmTjN��.���4W�0$������j�ܔ�Y;b\!�z��H*@1�p�*J��l�ʌY�^�m�J���J�u&��������߉$Z�rz�Q�B}�����)��i���Vn���te<�h���+��~���
���t^O�#���7��kH�����~̍�_'��3;�ڄ�?N��ʹ8��CeJ�^Ϲ߬=j��i&׵0��
3�+�+@`�63�����NyHw�k���nmk&-��D"t�ђ�� �@����0!C:�^��~��J�KP���w��1�k}�[.��10��PX#ǉ�=z&����Q�L���'o�T��a0����:�i��\Vʆϸ��0s�Z<�u�S���|6���_���I�pWk�$+`�ͯ1�#1?]~��BA@�F9O	�q s����࿬8?����Ӱ.��T�:$��NL3�w��e������� �Ǚߺ������1��l�ؑz�ws��N3�<Mhw~��{Q��LSI���B���j�d$xd�_�̉{�>�$�5�3-���uK2/zQޠ�z��(��ϏC��B�	�� ��*KhT�Z���mf&��}�����x%		c�C�F� N�O��*��#{Gќ��uTecpfb��_v|��fpK�����.u�Ht���M�ī>�q��a���6	��jA��~�-?���A�,�]Yt73����K-Jz`��{�c�rJԚ!�m;K3wD�<*�z�&ޔ��[g��&�Imc�yٝ��qw�ʟ�����J ��Φ��p�U݌^���U�v�Z[o�g�I
�����k�����X�1�v�/~�K��n���l�t���`��Y
ث �p BN���%�P���ߵ?�U+ ��������ȅ�߶_�X������$��\
Z��~0��A�Z�s�"�0^jߓ��L���])�GV�P�;b�\�c�~�^^P���u����q��Z�D����3&���=v`}.�i��B�&�U\P�3V�~�i�QU�*r����hV}c~#��Zw��k%i��k�.�#�t�[�^2�p6n�S|zr%��;����rA�f�`�+`�Lz. (.�Hfr��~�6Iy����jAVǒ�Li�CN��.ߛr@w�
�Uϴ���9>@�-����׆nVO� +;���LwP�0d{���ܡ;}�]�zb-�$�^ۡƊ�����-�?J=�YB8�BЁltF�Et�G��j�v��^�I��%lĉR�-6��K��󛑸q�z!��!ֈ��t�	X@>E�i8��kGg�Ɵ_G�Z�].`�q�M�1���F��>�~�jކ�6��=ܟ�f'�޶�WN�&��2�� Rޒv&��u�L]NB���e]p�J7�_J�`��]o�.vB5^�W=,�w'�z�Ten�Z�Cȧm=[��o뙟�}q6�n���E�Xԛ����Wcz���5�÷|3�qj��G�R�K��k�^�	�|�.Nk�K'	�Q=v�t�42�X�*~մ��gz?ߞ�q����TH\E�R6�DH�h[�ϧ.o����(�&�|���b��ǡ�t��P#�{�1�5ް�\���K�� z>�+����K�h���] S#v�Q4�I��bv��"��Ɇ�O�ë�_H�::� �q+$�!�Mh�WW�c��mh�TD�J��|PG���u�~N��w��Z����ڜ��S��"�y<�'��y=SSdrUʅs�1�4��5����8;����-u��HSAt�eU��՝��j���Zk�>\\�X�Qؤх�����Av��-@�!糳�Y���+N���S$1�e\W�W�%��"/�^�����+Q��Ҙ.P�Z��#�e�iUv�B���I�V�
�#�(鸃���.r����{�Ws�ɗ"��ݡ3� ���43��t!��֦S�z㮵���/`�9�&>���C�;��@o/�!��n�[�6)Wm*+�,̷488a�[e����O������|�XD��mw�s�VI�ʜ�e�����m��#�U�֒0��1@����`)�vW��s�i{�n'� �s�Z�����oR�W2k���J�,̐9��x��^�N7�͆�o�@���oug���m�����I�}kռt������>�֬��[��A�R���K����0��{ȏ�w��UK9D�&�+Ҏ.�*o��c��u˶�zT������0Plz�"l�C\�|��Zb��U�z�p�qIR���ŵ��i i����@՜���n��8~���닰��N�y1wW�r��P��9��Z#�U#y�L�Y���޻������V)�����G�L>q℗K�_���Q��gHF��,��Џ�ԭ�=ϦE�����`�����������_�
����:|��r�sw+/�\�l�+��9��7�3okp
|+L_�t'�����]�Q�����ɾ5TK*L�
�]U V�:F�^7�CV��a���$V�6��s�g`��q.ě+0
ś��*R�\������z�Qj^���;'��+v)�8򵐼�s(��E��������'���ʕ~Wa�����]#7s�t�me�4D@�����WY�6��2������>��CB�S�/�e����B��ۑ��;&����n��x�ݏg�/]I�	�#;�ӡ�JO@6�Xi\0��:@�N�7�Cyzc�1��n4�8友�J��O	��-Ox[C0��=!��cj����e|s}v-��M�`I)W&R���p���gחr��g���v��y4}o��T�GP���HQX8�FK��^�~��Obk�J>#�aM�y!���Z�A�,!�N�F>�Dg�;�8��e���=]��J�-���ϊ��<#�Ꮎ��r~:�������2n�e"��x}%2ʶ(%�-�?����V�����9�׳�s��\3.�po�u7��s�v�Y���8��fN	�n:�=s����4��l��F�!p|�J/���7f�y���h5Т���p(���{j<ͫ����PNRvt���@
7W~Q����2���$b���J����k 퍕���вd���_Y��V����x�X�Ulڍ(e�w͗?�3�&(�3�%9��?�}�|�E�2S��K�X�nX�C�`� 	~�'}d�N7օxz�~�n���b鄹]�S��*��e���'=�����u�-��.o6�fx՗F( �Fz��(FC�'��Oq3?�����} �Ӡ�6��"�+�/���ç��ѧ.YLLR�^hxD��D}��Ԙ��@9x_?���7�p|�ȋ����fUJ%.X���]N@O�F�.-y�E��Z�2��ʞ�-��N���Z��xh�����(vx-�7�9V�FM�>�!O�|�^�� :;o�S��-��A�O�L�~/Y﴿_�XO��YL;�^G�� ������LuJ T`K�3	P��C���OSL(˫��Mq� �0���>��4�2f����Y�)@�}-��g�+�X�(6q�u���8�*�z�
�"��n�0χM��*`��6�z1���>����ƿ��q���)s��U�2�f1���pO�d$�����<�3�2%���A쌑GX� �_X���4wk��@_�홐?H%�hfu�!�v��p�l6T���[ �z�_��}'�R/���@�[�ݹ�{�����?B�� 5�.����Kے��`��㋣׏!����24�wr#�~J^t5��R��_+}[l��]u�,����c�L�G|�޽$kB�vg�|>�K�2�G�Ӝ�+b9^U��nk:��T���C+��.����Y�O?OZt���2��v[������ ݷ^߸K��['�)ֺ�*&�����)6M�Y=#� /2��Z#}M��GU�.��F�>Y�l��-]�y"�1�y������.3�Ȱ�^@�<�>���P�r��(���V�j60���a�{:Lu�'h�~r~/�$]3���M�m+0��ڂb�M�*]�����e��bQq�8o�� �z��q�޼jy1+�Y��/��S1�N����+,T(�Nki����~��n��uIx~�q�����>�**��f�ވ�d~S7��ï�#���n���%]�۔3mAya��#�33��,��P�%,WId��E)���	���S�a�6k��=�E+~���Іgyٶئ3x�ئ��'���n�1��d��"p����v.0���x���`�����(����FYF`s)^i�P���F�(I{!%`b�W��7`�"e���L#�>�S9DI���e�,��o����p�.�*|�+a�9q��:itSd>Aϥ�Γ�2�Y|��M��<����ݥ�\*ڧ�cl_��?	�����Y.�������^o?6�M�W�"A��>��v�+�W\>#vV���=aY����^�xy&:�:s��F�wDE�Kӡ1���wl���U�9j��GaG���_H����2�p�F�q��ۅ���|N�1;+��o*��#]6��A��B���^3������M1�<��%{���f�^��������ٛG��M����(���6�=;��'�;t��9H�c�o���K�w��\���.K����d��j��jU3����v �"�4AF��;:�;�\�s�1��� ��O4�T4�`��F�V�\�և�ZUz2��o��l�	��0u���ei��I���b�;�Wgk��n�3%ϷW����ߌ9܂%�ދ�d�+���no��r� ���K����^O��=�ɲ&�؜ry�`�o���I��w_)��u6���}z{7�Q�s�1�����������n�ă|���0��D�+d]Z���A��er�Cg�����lֺ�Eb��˙�ms
�.�:���g.z�<պhG�����eG7hxv������I�+݇���O��Aj���$\��'O�3��"|��S�3_�vk��۝7m���Q�r x�o@����k���ޞ�x��s�����,�2��NzF�~�t�~t��j���M,�}���X�ӜX;�|t������~�(�^�`lA�
+�����"^�\��5"���F���E:j��X�s]]�띥���؉暑��7"F���!7~��L�;�m�K�1�)�K�\�T��*Y{��\��G�(>�Th*�#={���`t�j�=s�ڋ�%��4�d)�h���u9�o�Y<�3<F �1u)���1����>�;֕66 �	�V;�H#9�ڸq�v��Z[զC��JL�%�Ua{lI��w�20~��NOO;��̖���.}T�T`�>s�Ve�+��ɳ�.4IǗ��ߘ��mй�M�Ð�"j2"�[�jHȁ���9,υT���iE�7v�X�}EC�V,����B�.=��������#p�0�)��4��k;�vi�C@����|���o��}}o�%HY�0���xLp�n��̰���Έ���ȭ��CmF��q"�R*pp��p��`�r�Ή���*@K�?��[�����fk��r�����1Y�^�.�+�)�A���g��J����܀�+{�!��r[�?O"���mg�cL�Z�d{EW_�`�{�Y�͝�z��,-��wgd�D�!�o��9�I�9kOV���?��C�h�G��}�Az��QDK���]O�h0 }�S�Jc�V~;�!I�]�y  ��_��ʼ����@�����7���(`�Q��ɭ��PDa	c���Q�"��c-Wi����k�s�b�ؘ7�Ŧ�W^U/���qM�	�2$���9/��v%}7�����<��N���)#5��;��,��o���-�����~2#��I��c���"-�MNp{9���k�ZG&�3瘩�Up��؊�F �.�o��U�ŵ8º�,�*�|�ڱ���a-_��t|3_�ð�J%���%�����7_�J%�ta|[3~�h+;O�9YmVl�w��|������H�P!�oF��9J ]ٷ?��vU8?��'����Z��N!I�e*,�e4 B���ʤ��|��g!�6�t��=�RO'E���z�w�:6�B�b����@�Fg��tmR������u7����P��[t"W	q�u%݄PCNd�8O~.���d�I�Qb4û��b7^��&��t<4��24��Id�]I���<�;�&�l~5<�G�Xj��{�f��QLV�(�C�me�_�۩�و�ȯ_p�[X�Y����y�K��A�P�;�����%وhwu�Ne%:�[n�����A|�B��`���{�?���y�T�`[@*�j5�]�w��������`��Q猹�����ob�,jEW�hL��ĠoԨj/��Őj硎���j�4]�T��Ydv�z�E*CLaZan�Z��<;I�*]�%hL���;F��|�"l�����BK{{�Ո�8�hȟt�iQ���\��k�'}����R������̏1�R��5c�#3����C�{�GZNX߫A��y�Yĝ��*�µ��҇\)��{F'S;��Ck�GE\�e)ӵM����!IT�Ӆ1��̺c���3�m�y��
�<xk��P�~��?
�̜aV?�'f���Z
�1��7�Eg��('dr�g�&�p���`���/%�J���C.�	�5���D-L޵�op�?�EC�͕E��[��t��m'�7�T4�u���)����'�d&�Wv�ں�ԮP�zĕ.R`X��V��-~�d�C����3EbWi$C8(:O�5~��O�K-�p͏�J���f��]/{�
ʶ�h`�(����"~V<C�]A�cre��Te��"-���
�G,��̸H�2�m�z��P�<���DLT��W�nZ+�%�(�IP�%�FA�aH� ��V(�T�:�#QS-9����B��s��5����z<����4�@j���lL����-��8N��L҃*jȎ�$ *��3I�ɃW�ޠ>'u_;<�!�K�I�j�.�>E{"����Wp��u�ցR�Kqw� ��;w���R܋C�(�N��� ����\z����1���kMYk?9<�G��i��)i�3�m%_�l�������g༈*Q�[��³�O)��R/B�&���3;��`|?W`�>��>~���ō��L���oܞ�+��N1�D��[i������8�S��x[f�Xc�i���W�͗��`�G>���Rj�QJ����.�^�<`'�����Kj�r�|'&������5m$DA y^�x+2�J�ʚ�(�5�r#�� s��P��R�b�WGܽ�a�����ߪB��Bu�R+��o��
TZm|�eC2���l�T<�r�b�xlU��-�����&�b�����R�b�ҔF���}�~�k0���`���0����l�-�}�>��l{4�*M	D�i������nUx\
߲�\�=I'e��A2}�{�a���@وlˏH���f��e�$*1����A���܃�[��zi��,��3�Hލ$��X�ܯ"�鿯�)�/a�|��rH���,Ɓ�?��K�k��יO:�?r�-���L+�NGݚ���W���,"��1&�	ω�O�q�ZPM�`g�R����3yV�E�la�O�T���I�a��6�ҟ��e�ߦ4�>�	~�/O���l>T~j��D*�C��T�5�4��V�Z��;��|�>IY�;�q���Ç|î��ϜC���WI�i���x����J�}���i|�{�V�T]��'C���s���l��+�<�Wd
��<��=�%Τ6>b�酁)���g�C��Ul�JC!n�$([	x|sh:!��j!}	v��"g�T�΅�i�B̍O�2ظ��]�M铘��EX�'dڂ��!�ʣ���l�g�m�1&����^p�M��#���v5;јfڠ�tR��a�'��u�ģ--5�U��_�]�,m��<SZ��"�vx
��uj5�qWM[�f�c�zt��\ۭR���/�c�3wN�_4 �u��ōo��_S^`/{^�4mUb�y��.��Y���d��ڙv�<���e�e+��f�M���
�2O$j��/�_,�����q�N3�N6�?��/o��+RO�d)Er�y����2���_���3���gv�+;��y�����]y��	ח���6f|��j6�$�o��K�Dt̜,=��Y[�+��K�IG���J�rJ�w�(z�c�b�\���Sۍul�J���R,����ns�ӻr\#���jP�6"��|��}���&���veYY �6�!B��I���ڻ	��f��3[��kR�W������ɖ��D�㘈<2f�1�c~�6֩%�ݺ̜_N�ƻ�s�lE_���Y������:�T���m���.s�ki�m��U��� ��v�*��3�r��>c�D|:��� հ³)Kuѷ,�4h�5�/�L>{
wC�����ޣe���D<�ށCG�S��9������o]���:�ƙ��MPS�%�ca�{z
�x��*����3o����
���[&��!��	K
�MCH��rK���@iu?=������ۿ�-t��L�+��F��Աz�՛�����A�wG�ʳ����k�E��ޔX��R�����Tx"O�s�����O�6T���8���vaOU���0t{��I8N�	�g��6셔�����y��|P�ۢ�j�zQ��f4O��rlh�v��ʃ-�����嫧魊�{Ζ��b�K�����/e��&��v*���;�6S�Y��7jk.ϸ]2�x�I�?7)~�I;#!y	rx@�|*�?~���Tc��
,��F9���/	�c,+T�uW���B��l��U�����k�Z&��TtN �^Ó���E;'ص�z�r68��,4�	�R�x��x&&x�0|;h1���/���w��1��bH�P��o�x����̋#"�db�Y����>�V;��c��>���W�ţk�Ä9}����ƣulC�}����Փy�$��Y����^wVFc�bHt��F��󦂌����f����^�\�$e��G/P�Oid�H�9Z��ڙ�'H `����"e7`���'�
��
/}����e���8�^f���br��e�?�������2y]c��x�PS�7>�Pi(�W%,�PG����R��.�lq����D�	�}5.K�� C��=c��>��ll �t)ܙ�`�k�`���	�U�B����I�y���)v�G���v�ǝ:vV�M��H�ú��!  xU�������
˙����Ej�"&���n=�RR�zLMmѷ9�<�P�PV��
*�8��B#c�\Z^�>o�Uޗ�J<g%x*|��P.&��:��=n�V�v���S��%o��o�7��٧*��С����!n99�a�t�,76-�&�o0�R��l���&d���|�T���������N�Xﱭ�{c��9���A��؃�k��ʙ���X�j�Izoc�^s5$�V0f�׋���:�+��sޢ��X�e�[#w�m(Lv��Z�|�}�/�Da�'9�a���ѭ�ˀˌ�Kd�H@�ޡk
��,)�t�J;�O�#$��%�<�8DJTk��Y�����#�:���Պ`���5Cս9��V�稔])l.�����=x�6��%v�Kְ�8��۟q�7�b6EX�p�|s�� K���ߣd�qOJ��_�Bd��_�����C�u�X�/2V�|�V?n�r��;P�]�Q�TVI3��-���)�o�+����o`� �.�����f3�y!��3�XBқ�W]�]���i�����_���/эB�qY�~����[�dڠҎ�A�9���tK��hls�������������?�ō������!���*��y\�C����q���=,�����66B����M��$��7��:��9MOf��JV^n5�R����æ���MX�A�v�#ں��k6�z�/�f�bZ#���AU���)L�j��s~b�)����v�z��x�Y�h�������&�ٱ�;u�����$�'	;�-�-�n��Ɖ����
Y�Z��׍#�u���}ɇ��Ly��ɱ�@���M���̋��YCk�qca��������qQ��
r��D�x�CY�%�V�_.��[5
�Z��<eB!����O4�g�����Ű�� ���
]�x�Fs~��u~��)��B�-f��Ձ�ƿ
q�?0��7��MW�����'�x�'�کň�.���Z^=�d@�_�>#1ԉq���%+�� o�1���n�S��`&^4��A���G��w�J
�>s�CWn��ԁ���σ��b���(��a�uNf��R�s�[�-��،Mѥ^0%�%�8Ǔ�\��ϻ�<Zˁj�~�c{��Nes�N��ϲ6�n٘���ZV��&����E�Qnb�N�&�ao[�ӂ�+@����*�l��E f;���Fz�	���@>ĲI��Wؔե5��f�3����	����1�ê���ʛL:L�2"��r���
\�K�3י^�^$XU�,���Ef�z�'�Ҩ�A��~&g�5Z���i��QI,�ߩJB�O������1F-�Y���}��w�l5[
����p$�M@{�p�&(-���[_�Z�:##\�SV.َr�?اfӴ5C#,�磴��ԛ0��ͱ?v���D$<��nost��RO% jSA������dy���>ȝv�*+)�(®��.r4|�2I�󧘈z���	����2���Ջ���A�U"l'���"���~ǐ���,�d��SA�:
���\sl�Q�`�D�����)��Lv9|W�p/���>���h6o�����,P^������4O5;���l�{�߰%��bm�sW/W�ה����y������]ZU8S��	�g;��) �=���[���1�df���XI��A�X�y��[������>����2ݛ��S�6	�pB������D>�Z�I,�5�~��L�F�#�xш{�^��"�k���z��.6�a�������!�1Tռ�(��y�b:�-k���E�4e_#r��;��-�r"jM8�Hۑ~?)�@����}=F��g�p�y])�-��ɼ���''8$=��W�cDC�Ѕ�2�۽�m�&&��w��-LPC�a�d���O�&���1W���ʝ2P�VoK�Z.�\��"���!�Co0D(�Q�o��� �)~��H�b-,��U���9؃lK�V��}�/I�b�4j`�jL:��Gnt�E	��Mߊ��mA�K�K�+�2����&����CJ�s��w[����[Q-ȂB�.Qi;?��Z�(���sJ�F��KR�̏{d�}V�����#�y٥#x��n�q�,�hzC���xn=Jc|1a�AR}�Nߴȍ�zv�O�6���>���.�7J�@c'��N��>w&x���[�7�\��GQÒ��|�zĂ�/�c��\N������Xu���7�����T����!� �}�N�'�r�g�W�z�.=��d��D�(}m�Zh�x�k��>e<=0�5��U�uIZ,������:������Ki��S���I�Ȋ`Y��p�~��%�.^?����T��]�,�����[�G�Fw&���j�5Dng��S��J���V�����+�5�i.��!̂Ѡ��V Z�yO����j�Q��pZV��(+1�g�|�+�OϑM�N&�5�/�w�;/�s�c )�t�6��'���O��ח
��ٮ�%O�?�τ$��J"�㦅�BQ��;�`q� �0oEU_��YM�z%�#�s�o�-^�@f���v�6?;���IަGJ�iG���Mo��Tu���r	��ݝ�v��ְNK�O��,�Cm	^n=��D
~�<����w�W���\Dtp�6¨��r�i[�{9�*��z�eaf9�=:�c���t�WR岞��[P��z��
WIzqi��#���C�̥I
����|6Œ1�(��!�ޭ۵������W�C�����Կ�tm�?��j����Nĩ�]�x:9��mO�<>��jS��V����2�T\�nC�TG�`�}+�7ʉ�,�^(��nI����H+�/�	I�����%��0�cȿ�h&�M�`'����wLUS�ő���ڂ����R�5�]�mk����<�OA{��'�f��e"N���v�(���ͮdT+2+@~���
�k�ժH����;�}��C�;3�_����2����Pa���/DI�N��!��f���43���������DaZ����[��F ���
�?8[��/��q�|j�V�^���X(��r�S����K�$��r�`�dVL#�!�0���2�DFKO_��0��/�a�x�X���R�f�m�/�_.��f*�-���oԳ@1φ�I.53;=3����y���-7\|�pr��+�=+���l���|S.lcƠGa� ��@16V�0C�6	g{���c�8���1��~{d�L�[8����T�fl��O�̈́A2]�Kz�{%$,JMz�p�PW䉴<�5님������;ZO��	�p��rx�/21�F�=�9��t�e�yr�h���yO���}��V��>c仞�-,;�7NhEO<+�fUyU����i�͢�ߙ�6^��jΦB�~�z�O5�:�k�m��̴�e��5"��ѐH0n�4�Z������[��σ'`��(1�ɟLR�Q��aW��g��g^�F���B�*>��ŦW�
�a�G�z��$Mٝ8v��Z�^�8��6"l<|���Y-ەb<�`�[��\���u6�ny,��TA�W1�Y,�o�w1��>�w�y���"<YL��T������ �J�#�kC��O�n�>!`lqf2m�z�Pb�r�mf��ݒ�x+��5�`PJ����Z����gh�X)ڌuye��ȣ��c���.
�Q���u2�RHV��k�2;ү�lr�A���ɷ�n%��䋿tt*!Ie�6���ws�e������v��j�O!��9�L���"V��K��1~��H��	o�������?�_��2�V��hƛʘF%���J�W��D�1�Y�Y��$��F���x�DP��,[&x&k���׳����_�cօ���H���.��a

@�S)�h゜�A�~範I	Le��� ��a��S���"8������S�Bo␅�@?�����s�:�w?�.*V<����i�6��s{9T��b��wqU���5o�h���q$�v��Х;mV�S���N��:�E�۾�?�x2�=	���Ebڗ ���W7����B��4��n���t� '��(a<�Fz��Z�%�D�z��o�x��@O��ZU����gļ�tw�E��v�^�>2����	ARcU�G0�n�p-dcPz��M)��g�c����	�wG.j��f���.F�o�Fb.$11l�$-��f�$12�H�:�f0�	K����ޝY?8��P�X��ԌZٶ#�U����;l�mC�z��I�݉[��|��J�d��qK��p��%(J���p�S���/'��#�3)7����֥������v�^o�TqhD�����wJ|l|�6����qUS�Cݦ�3a���>��J��|hm��c���Da��u�/�<�zk��Sf�]�I�պ,����;B�욌�R��E�1�-�� ������h�}��Ej�����H+8dmow��-�$rs����!� �mA$:�`�0+Z؋[�|��� �H[�ئƚD�Kg:�>�
O��-�n��(�Ѓ;d�7��*�����~��r�^�"9Ɵ �w��G�4�� �G��&�:w�:="��c�<@s�5�/�o�ot"��7��c:�r���X�oW�����hf)�?�P������yJ�L�@�q<Y��m��R�����6,�r��1Շ����?�Q��6�4�f[(��u�lhR�����`y�h��(;�=��b,
�.v�u>]�a��t��ٝò�|�hN��s��n��Ds��%�ێ�(�\B{f~��wP�;O]�q�e:��|:��ñaX�<�jfJ�!�ߪʝ�&�#�~q�QA���nT͝�ݻt�7$���(��3��꥖��GM?
��@QR�_�2��g17�͑aR�SB��0�"S�r��_��oP8-�p�u�{K���^�_��䕄M~MCCH�$8f�]c���n�;yɑB��{���.�����b\�Y{c��`h���	���<['��t������V[h�����Fhpu�AҾ�O,��������Xt��K��O���1D
*���6@q��^9{W��xd�`�B��5�fݬ����D�N)�$:�,,j:�����C���w-2|K�J	�(��yA!���WS��NV+l�5 �$H��'�(�c���_L�~��~�JF~�����m"x�vw�������(2qW���F�U��8b�+80^e̼�Z��c�c��J{�$҃o���[82�y6�8��\�f)�ѝ�恎�wK���=������^�형�ƚ���}8z{Qw�阀��A�|��nj��O^�b��[��l����i����#�@uAS��v�lk܍ƌ��RY�iS%�@����7�:�nH�jxO�q"3	�h�-r��h� �H'گ��=�C��o�H���^57cb��p��(��Fٻ`꿃G����_W�(M��~�U����2ic�ǖҖ�}|�+��E�~��[7�?��Ǻ�����a������!�)���w��}�����m�����!G֯�>�v%}�|�H���A���Ͽ�+�S�X�M�/���H,7;�p��.D�G���=��q�W|u_�L �r=1
?�b�-s��8?�;�k"Ra��D�)~�F�F��N26+���=�K�6Y��E�w��+����k�D\9���N���`?|l�k����)�����O����S�:RUO�=�N�]K�0�����@Y��y!�J쵱��������%�ٍ�9WA�*x���R�����R��[6νmϨ�K�� ���m>��w��˧p0��t��4t����tۭ*(�͢����O��� վjs� \���lP8]�!]�c	/4���j��X�6V�7�YYPOC�b6�M���b��h��. $}B^@!�Kv�g�d�X~���`�}q��!���z�NE&紦�ad Ҍ�z�Rd�Щ�������3�%�Y��\�>�4�z��NP��D�-�x���$���ͿZ5*� k$����b^Tբݔ�P^�x+�nt�߄>$��g�k��0.��q^�.�Xi����)��VQ��3ܩmV��"�)�D;���3�O�/z T�ن9�5{Ĩ0�V�M��C7�ZA4x���T���Gh���2feb�or
�p����G��|�Y��j[&8K���_1��	�RG����\*7�+b����e~4yqud�HZ4������a��$���=R��֧���l��*�6٤Q�#���e��Y��~�-��Emn�I��'!摾%*V��w���	�4F�Ҹn��r���	D�o1~��PeB�?.H� �<3����h��?�Gy���K~�����u��'�U�n����'+�[���c^�k[7U����Ǜ�>�BH�Q��b(�~ +����k��y�t�[=�.�Coˣ�t]�"��F}@NF=����T�� d�9f7������4���ףb��'9�Qt�8:RgE���KEUn����lϫ���=JkH L��7��d���>��)�t�y�<~����e��R���曾ֆ�3��&�,�_]W����	m��%=/}!�aZ_�s�~�xs�
I���gj!�5�+���<��Y�<i1���=�Q9K��"gD�6�mS�%Rh��q�ӧV�@�-�^�w�"Z����G?��<�j� Y_71^�1� lM��]R��I�+��/V�#Q�١�YB�����_�ں����<k���ũ�11=��� �*pO�t�ů��N�?�+Kl��j�>��x��#�qm8�_YQ3�ӻ?�m�,%v�0JN�����B����(����^㆒�>ip6��+o%u����֣��3�]���|j�������&�1]�F0�UϞ�|��I�[刦^�]鑢�fEt�W���e���Rq�^�T�w ���P6�z`�e��N=&��/��5�z�?Y	��j�_~ ��2�W�r�⏱��鵔���G"��a�|���B(��G�})�Vъ�!k�B�M��/�'%i�[tޱ��ݵ��T��;u�/|�y���\��Y��{��0d�%���fL������Vd���m�;H�E������$�q��W�'%�ua����ĥ͎W�Ǚ��~\��o��U�Ͻ�2Г[᪞���~��s�S{�2G#��WGǷ�;��|UY���&D�S�g"���&:/Z`!�(ף�Cn<��{S�J�b�w~�����!�4��:ʱ��!Z�[�ِ�m>����ͫ�A����QL��X�����R��m�^g�s��;��3c�v�C��{O��$�X�H�Ť�f^y-�ϦV�;�E���Z5�2����"��Ī��f뚢|�r���W ��L����6υC�l�"�?��6CN��Hl��[��e�����ٿ�<��xMeR�C�����Fѿ�n�C�:p�����Q�+
��eT,�?�f�&�������O/>.۫��Sc�����a6=s+Z�o;׶�p�b��Ѽ��Mv��`~S�=@*��-�bͷ"� �~m=[sW�g�n|4O�B�����h�1fmQ�P�U�á�L� ���F�]�l��yt����I��yQ�qk!�j�7�Gf�S�]���B��V� 9�b`��x��QH�[�^9�1��gw���%6H�z"���Sf�w�q����o˙>��H���Z�i���<�0��w��<	9���+���,L=����N=>3���2�!���+Mչ1�3� �F����L�~��^:g7YWS[�S�{S��_��oߎ]��^B$v ={����Y�gz®���ql"?vz�	U��"��.��K�2D�E'�'~+.�Z9���gט�wI��D{�v�L�QM� G�viŅoh�����k�S��֝]�8	OAWܖ_7��Ki����6i��5��Cb��-Ò����s��Y"}�pT�6O_ U�.`E�K*/y��^8���/0��y�L؍�)E����~gI����T�ޝ|=�mM?��X �<�]�����+>����Σ�8�mDMs��$�n^�����"t����o�6�v0��9�o���r_�17�����گ�QwG9��-
�:M����a���chGM�m�Φa ����⺃r,3���^zH��?ߠF�]��ax�j�s�2^C`d��u݆~A#}�{��V�Di��}@ �D����s��uފV��@����,~���r�l��*)��������T!ƅK�7:�o��nq��i�����,�P����}�!��\\X����R"��Wg�R#!1}X��������@6|A��d�ݬ�����{�b�M;Ь�h�n�tϤm�=��ӛ���Q/�5۾P�0��_T��P����5�.��J����b���xt>MM���6�-	��i����?����qT�(���3�渊.7�:�5���eo|��f\vMq�i�:�3��vz���Q��Tz5ch�/�0�t��7$��Q��������g�+r>"Y��8��Te.%;�7�
��߉���ڮ����؊��׼��쯺`R2�U_�3��O]�:?����*����/��HS�h�'6luf�P�	�@�Md�I�t��\��WZ/Z1#<0�]�_�6�P�j�J�Br�����كP#����is�#�I%��sD��1\���U����� ��SS={�_C�3�J�7���	0>�L�e)�U�j�b9�?���]��"4�顃Kv#'�4а�wl	�aO�J�L,�<�E�u�n���޽-�����Yq�&"(a��t�8��n]�'h�����0	��٣*�Me�j��]�(kEP�/o�F�6�t�(��<Y:���EWv�ޤ����t��$;pӦW���x\�'\	r�&���nN���w%�{wG�S��v\)f����x?;p�e瀲;�.%�f����t:�@x�q�r�:�a=6���2x��v�%*���ʎ!e�]�tM׼yn��.y��)�M\"7�rC4�-
�v��筥�C�V@�ge����X�m~�D��;�m��bG���`6��A����Ҫ�zO��̛��P��.^h��<�Y�_c�Ux�d��3�?��j����b�Mf�h�)��W�v���>4f�S�z�6M���֢��i�̔�7�vj�#_��կ�_
}�4 ������\�~���#����5��ýz��p�!��u��Vo|����[�h��Kb���^�̡.l(�`f���t���O�x9]K�^}��h�B8{���95��nߛ�߇���\��Ů_����A�'s}Ju����X{�qtF�����jUh�r�;6�o�	E�ڤD��#[/7�\��r6��ϻ��<�9�(��i��-'�!�x��L��S�h�!.���6u���N��3*-�X�O�]Hz�������KX��Rb	g���i������z��#�Wm�k�;��-��0 �L�������z"�|�}�ɀx4��Fu�5'��ʋ���MҤ�Y��љ������6f���|YF��A�[7�щ�#ӑ���^�����9o^�6E��zA"�D�U3�;�f���ؚ�T#�c.Uמ%K����VʀAH�J��^D�X�!�����mK��d��G��ݜ��`�$���\T�ǅ�N�o?��j57]z\{������j�8�$�� ײV9��Ѫj���@z�ht�����ݬ�Ӄ���һ�n�-{)�w����������5��Vܧ���0�&�f��Ԥ:�I�Z�Ë�3b��8x<E9+E!Q�[=���1فl�+�20Ə��7�Z����[�tϛ/n�8���X���Пl�S���6��Ӳ M	�H/:���z|��PB�aMb&���
��v�δMK_�h�nkJZ����6��� )���]hד�Ǝv y�K�*Bq�l��mRT�!s$i)�M����e��Y}~[�H*ߠÏ��d ��ޏr�7y�6
rO�"�F����2���,�����C�n�v�� X�U�ڞ%V����A(�*�=z��"����(%�rx�_)�������lNU2�f����WBd�'�r5�x����@�b�6��4q����o�4�R���������>]o����+$H�r��?oH���ϡvPK�5o/�S�=��u�[�Mf[�R�/p��)�v�@"�|7�**�#�B��8ţ�wh���ՙ��]�G�����(��]t)�I���ln��+�;mS ]6a����5��]Ҧ��ͣT,E�et~ɇ{�/�drW�6�����|hymR��G�\�B?�x4�B�>�2�'L���&~�KҴ��tV��<�J6i��b:��'O�����m8ylA%��<;����J$�����&1��PD�P|��}�&F��F0�E�\w������b�Ae�:��o!Ӥ��-��h�$F����a��I�����K�^p��� �b�\�r�O��6z���g�&�K6���<����q�m�ǽ4�Y�ލ��M�]�.��\gQ��yֆ�%5�^k�"u��)aS-鵳K��*�ϟ	���r�{�e�>BL��k����E9���6�^o����Ҟ���yb���Qe��A]���*'���i�0=�@���R��	{���G݃�����j8*�^��������{&��%�6_�\��n+�Y���9�򺯒g������eo�>�*����f(��`i�<k�AΜ����Q~o[�0��=���ۧ�<u�n��m��~��#Y�PWL�nD��7�}p%����j���ȇ������s�_�"i�fr<��[��Zty<^��~Pd6�ߴ�h��2{�ȏ����Q
!����GO���E�h:m��S��V\�d�n�i9Ϙ�������맘�~�z ��Օ��A&@�`J�	UϘ{�B;U7�ڬ����K"ot�m�rtm�&m �g)�3si�[ep{��%��:���6�ݠ��'Ꭰ\8d����;�������6��df�V�섩�c59Y(��,�8�Z�н#��ӧ�2�1� ��l���gl2�����A�s2����嚤kX�Y����0�:=?Kc5��2��T<��{!f���{�'��ޕ�����}BtR�{\a�w^����&��W����%B���^u�͓���8��i�;
�U�	���8�p0�`�d�Ɇ�}c��$v��"��I�p�:�]��<RE��j�u%�f�%h���Q�]t�l{;8��q�݉^D�R	��Gw�mB��]�L����jpЛm�O8���K�"���+cp�e-~���ag��W�=��_��	HިȒג2#w8'<����}&�m�連<`�ED:����&sg�">����^���.{�㚚�i��5"V$=B��"����N{����6�W������l����0�H�	��>(��W��b�Ju~6P4N�(,t���w5���w��+!p�cB�L��W��H����nw���=:8���t8˱a��@�l?>ἔ[��zڹɀ�n�L�G�����p�<BNƃ�"ۼ���8~����i���~D,66R��è
�B*��9K$�V}ّ�,�&鯗 :�kK~Q.3f�ӆ%��yK<���e����D�����Ň�\�?�b@;Z����.�[Fw�,�]�^bP6���Cj�,uI�$��o�;1Wv��4�3�S���|�k�5z�A�>U�Uiē7&�a<�����#v?/�q�G����7��xwO�n�[�M��ٴ��>�=o����2�ل�E2��u��W�U;��U�.G%��� ����i0��	IWVK2��Q�Ń�/��N�op��EPVŕ�̻�1�D��x	�lyg�$"yC�&u�K����������p_=�l|�@kA��!���p�D�t)]�)�Kv���̆Y��R���a��NZ2�Ê;��G���G{��k1���<ˉޓ";�� \J�߬�=�7�Nx�����2H���<)���=^����ϖ������O�S\�fU�:��L	G�e���#���{���\a��8W&�g���L������U�e|]7|�8 �$����[ڲ���D(&Rw��t��FN��f����v�ʗ�}����M�6��.�?�.��1���'��^�O�$N�"\�v����(�dpCO�ԯ���6�{�L�X$��W=@
G6��oRw/W�~���`�y;2�>h�h&+��0�l���RWJ;�R��X��`�04p}O�? 0l��S��Dߔ]K��n�k�b�\,ŝ�m�N����w���6�"�0#�$ٖY��1D�
Ǚ�V�0�?2R��04�����S�O�>��.�n�FsT B��33���.W�t{�[N^]�d�RF�|��\�:n_�]i�L7�Z�ٶ�Sl�*�w��hvPʇ�<��|7��s�\�?d�0������{��@�{aYsp�ba��.b�tr�C�+��"��~C3ÞnK3L�eo�b��pd�1��l�2;���T�����CI��/E�_�	tsF��8+�j�e%�}��ƃ�>��M_Q�y%�Ǿ�l2U���Rw��*rpjӻ��4�b�B$LS� &\�՟����N���}����f�jr�%��-Y-�{�c�Ę֮+��L�XCTi~ګ��+��_��9va��W\��G�A1�l�
N*�2_N&�:��#���w�����/�_���]��*W�E�h5�K�`��:���j�m�����dc�s̗�0+c�[�����]��ʥ��B@��|��m5��bp��A�F�K������~[�� ��N�K�d*�Ae:��ڠ�Z��l*��}�v����R5Zs�\a��]�v�K2����|�³!1���L�!���F]-7e��0��1-;�./���I��׉�T ?��]틕�7,>�d��4������9����Hv/m�h�%.x8oct |Z�%/�H(�-Oށ��D�:֝����.ZW��
.Mo��=�n�M�,d$��nwb_X"|
��:��=�����X`BhQy8	m��.�D*l��ˠ6Uc��I����uQ�m��+��M�|]x��!�cj�/E������AHR��6��������ແA�(s�NŐ T�s��U�]����^�i��4����m'��w��OV���A#���K�f�'T`���m�!��1��5-�<CY狤���)���W毿%����R7h�ViH�Hd�������L)Ju�D{���R MI`g5]��\A7�?����o�s���v��<�~_�[<��qи���_Nr+��;w ��߶u	%����ѴTZ�_�p�n`�Y�-�N�ն�{���dz��н,�d͐V��D�O�4��R�eU_� �����1�b���U�Eۤ	�!9�% }�������a��o��]��i�i^Z������Ǆ�yK�����P	�g�Y"C�{9d��^�GG8E!E��]�|,��Θ�$���ܒ@(A�N��y��X����QX8l2�?Qӿ���%bܳ�_9xqK��$������q�~��,���VʃU:���vnޱ�2�����Ӎ�y�q�g�*$ӽG���.�${F"nsO�"�D�_��$.A�/\w8p��!�\��A��
�1T J��m��	i�zτ��_�jG�}ݗ�|���-��Y������w-�;�.�g
y��S����a��HE�4~���_x�Y:e,_�"�د�c����Yf�ļ�m��inY�|T�m�����"�S\�;.��uŮ���zy�g��$���n��%���ʱ�}�z�-9����� ���Vk�kܔ��Gr=�?�)��-�pP�e$�����R�O�%j��(|��ޣY�@E�F�Ry;�Z]5�5p1�y�-����j�4n�v�?o��[�Xf�t;>������]��=u(���!�] ��ޮf�"��?��ծH�2kI-6[(�t�urNӺ)D�����v9�b0vLU��X��N9�T�;�@/��5Ț��G�����f7���29˿BD�ՀГ��6����I��n�U8l�x�6��Ye�ƬَE��w�G���\�>�%I�ߕ|�����e���5
;�<�����^j�ﳒr�៙�pڼ��.?ZB\H��5�,�I���)�u�J��l��6���ɽfR���r�Zb�� ��2V�)�΢�ͤj�Z濦�V�|�Ii�����y�2H�am~9ГT��j����:*�FJ�n6�9���P��[���O����
����� �#]�H)H	�-͐*��1�9 54#���9t� ~x�����9`����}��*SO���gYcU�w�$ݗí����gՆF�$K�)�eO��=�ϳ�+4TNPF��e�;�h�v�<'��(̳��|���e/�H�yJ�=?�牄Ξ͊s����fp[��(�\}�gWXK�y.�+UC����u���P��q�=b�ߣϴfH-�>#kni/o��"�!��$��g�+C�])��E�*��չ�T�R�K�������|�������h���[���r���b^��;��H�3+�e�a5K	���M�]�����K�'l�Nl�E�L�6>����.���֐����ШǾ@�C��'g�;F��u�^�i��+��
T 
m�WQ��SR��v��lB�2�=ШoP{�]5�]s�V��V�FW&mz;�<�Jް�կk�wG�p�ˑ�������α1�^���� cĩ_g'���l|�!��/�k���I�{K��Zv0�[��|Ǿ�;�FYV�|�E�� �⮒��N/s�2�]��6r�173e�b�̭&%6��:�
~r��b{T����ݢP����y��52Oڭ"�ʆSz�t�R�V u�w�yS\���*����nT�C�B��Dς��ԃ�L�k�Ȋ*���0/�䱧��]��>��_-�������?�u��"䐤%h�r��L雷r��;s�$E�ݍI�)P���,u���������o��M�)	��*NÆ[�)�/ַv�r����]�[�/�$x߇�N����<���h�hS�Ǘ"���41�|R�7������&P�/�a�g�z����7��_VF:����j�ƥ�i/�W`�+�r9���?�����_l<� �dR���Y��ȕ�`�v=U��=��/��:�S����9��Qbrja�ݠ����<ǢX�e���Z{o�Jo%�G�I�ͯ�Ԥ�ά�x�j��b&ƻ���|�a�y�Q�5 �_N�S��>w��L?9� �K�;�$���h����pI���?C����:�QA��N�ǿ����]�y�7�M���O-ɜ�w�&d�
��%5�x	�+��.b_�ZC�.�u����ʕ��
���gG{ڗGY�=����g-t���'���������+Eͺ/7)��/�MHt���c;*�!��t�ˮ�zmO?�f�����13?q%��Q�X��`��,�rY\��)h�}2���F�}:Y�Rݥ�gg��g�ۨ#`Peτ(brD.S,����w���1��܏��ؤ��ہdM�NGk��l�P9�Խ���-�ja���Y7s��6��e��V�G�v�����x�Uc�nDc���;���+j�E�U+Ͻ^�ˍ��7����'���L�qX�.��|r��1@�e��o(~���	�ߓQq@�ʈ.�L�5�p�~��,�3o��´�.���T��ଭ�X(C�Ң��[�¯�.�ݴ�;j3U&	�q
H�|���ڧH������veЭ���"��
�_7��̲&_^
 eK��F�OW}H0�[����2ۦ�%���!}�A\u3Z���Lb���B��-�z7���Iu�WJR�	���ax�
q��z�8q�~7TO�)��3s�84�X�ҫ�8�\y-^c��˯*n���l5Hn�&Ȗ\;Q���G%kl-�tG�&,���1�1����ͼĘE �`�ڼ &�4��M��)����Pk&�E�󜃦��=p����rϼNh�����9���!#���dE����$����V����X��;��_�]Јx(�\_O~I֋�qZ�]�L��*���X�R�~l\�(R�H�B!�d�)Q/�����cJŮ��k��q�z*�fN�IM�*�Ӣ����8\�l�lbz���X�����0��?J��u�&����E��=�L6
�|Q��'$9A�:P<�,1���/���7!��OZ&�-�΂�`�Z����<��ɚC�|�`�=/v��M޵�JHc�Y%9�Y� ������3Y�1��!)�#�h9���
�{�*,H:g�A���u	���ZY�g`��Ok�\��c�>�N��g5�Ѳ �0�.��s[��rW���"]��W�3����e���X񙮺"��CrIL{8�>q���[�P����k�߿l���K��+D����]T]	�eSm��g��J�u���`�1��I8��,y���T&Up���I�	�hm�G�^��Wfĝ`�JIe%��ð��X�}RBC5�x�D���=ӻ��}��<P�Y^����p-�W�f���3�����jJnv  ��f��h{���y���מ����<n����,(;���G���ۥ�O��ݩqIw)�=�NY%��c;�؋L{���Ky���f�� �5El=�9dR�B�&�A5rŀ�3غ^�۽~@a�ݻ��`�"s������xԌ;*��~�4@�)�G4�`�{�nC��M����'�2��0 XX��i����/4��c*�ڳi:A�,��f�ޖ����:��=\���D�ގ�w�kN^�x=��qq�1(���W��ѓ�V�4���y�s0�e�W�a�S���Xx+�y0uK�uu��w%�v�wӉ�Q߈�l�2׃;�?��+�8St��-����|��GTf�_�.�B}}y8E�طEm�U=�D8��2k��|/%6�{N�FM,ڱ�<a?&�24w�ٴ�������&��|4���8<��掕���
8|����K�8�;�.������!_wMm�&��c]0(3�(��y{�Ҵ�PPJ�.���Ş�F&�ր��<\X�R���Lbd��L�C*��/��\?������k$���Y�VHϿ�4Y�o$u�F��a��Dr�z]�2���*$�6+�UU[���_�B��U��9Lo��D'���_n9���[1Ðg1�� ���W�{e.m�+�����W�J���4c����O*0� 4�y�=���!�Xz����9��'Q��#�Z]W�ʏ�|�% (�Z=O�&f5k�����vO�_v�tZi(x뤫�_i�����9E=W��r8$���\ďg�ب�u�h���8��\�bS;��������&z_�����������l����ԯ�L�v�L?
�FUu]v�P���͒S�Q���(ǿQ!K�<�����g:|�ܓ(��F������ &��}꾘�	YD������X1�����p?�R��y�9��&�����'P����A����lۯܡZĚ$6%H�ƾ�<�nrn�Wӯ��la/�u��ݜQӄ����6��3ҎG֜�n��mԟ������ݣv+e�BvV��!��6�ė&)о��D'�S��AŌ��(�V�b�U�1P�(~p(IG:]�Qc��v����Y9���b���?�
e�﹯�
��	X#IQH����nVpx3��L�ԉ㺊��w���$�Z|* ���򭥒+4��d���I�ؙ�ȥ��M�Ji M�r����.��Gk=�q�ȕ�MN@�5��Tu~�I�+�e�SK�"���)6�*�P��Y���3�;J_�/$ A���j�H
s��Re���eV��F��F8A�q���yغ��ȵ,�#ŉ&Z���V�������h3�4��R'�v�Ϥ1zVޅ�0A����~�<$Ic�y�[���f�@��x6�8�|n�#�(�$`�f����\t��w�{/,�(���mE��bUXL�:W 򸴻J�+Sg�YH9Ʋdw�N���]M}������2L0E�^�;�
Y};�}�`d��Fl0�9K�x��,��L�gz�m,���nJb�F��]��)��{�B&��7
��+��k��.�x_��,���$^�5����@�����_m���/�t�)�?�U��iہ��U�L����$%�����
0)�
匹�=�؉��țٗ�su�)�˥ֹP���?*G���[���fzaԄ�4�BN���q��cp����=���|��%�e�Y(��"��M���s�ˊ�&.�#\�}ܻ � (�6�-z��;$2��������i�%���'�Y����|��f����n7��v3�����Vx��e��3��pӵ��_0��3,|��}?lg�z�>n�5��~z(~�����N�Z�q)��\r�\?vim��a�lN��E�H��Vn�܄;��:s���Y�֗{b?�\��z�q��<,KĭC�-��p�9{i�f�%y�<��ǡ;��]q.�1�[�M�q8\+-��7�p����ܴ�z�����(�`{�*,gx�
b}��|H�^�s�h�����I�z4<�}��f�8�ޞu���_6�Z8 ~�/DWY�W�[�Z/�ʥOJv�w���,$R|�K� �C����fe%EK^ָ%��؊5F�b �����qA�cARIH��eR >���-V�樏������</c�����u>��J
�>�v[C�_c�y��m�����L���Lo�;96�U�ҝ�@
���ϵ�!�hy�ÑϹv��gK>�>ы���vi3�*fX�m�Ng�А���xmj'�z�t�?_�ΞQt��7�w�������m=C^7��o�M:�@h!��^�བ�L-7�'��J딫����~K�
��*3�F%!Jٟ+<b_�$�ₐ�C��N n�i�����If��{���|��8T�&` ��k���M��er�U�;T���$��v��U-���c�Ǌ`��Y��|�ǦС��{��x�?���,��Q�MP��2�'?-�܏S�7nڶӨy����N�u�quoxe���XF;��!��������3,���W٢pܩT�tj9�E����gc(����QX-Fe��dm#D�#pҦC��,��>�l{EN=ն�P�ym۟�/�I\��Zzd�è�:Pw�U�{�ST*O����B@s��)�%+��CG��hy?~Y�-�K�v��~P��S�yϻ� ��y����M���y����빅�G���o^h��J�^ fn>�҈wh�.�}k�2����rQ�w9Cd.�=��e
i��#:�Τ���Y�'�Ӟ��>~2=սt��y�l�QWt��R@p��#��=_5�_O�F����^]�p�S��t�d�]���D������]��g���K�˝v���7�zx����X�w�.���U�L?)%�\|L����l�Y(�79��ž�սSq貄��6�F N���c��&��h&UD��r�s���W��6���ݾ�%�Л"�o���(�(�}�e=,U|r����b<�Q7 _�u���>l���B�	�;j3l�|"��@I��������l8r��<���_��E.����H����E�57u	<䀃.xe�*8IaG��G��߹�IR�u7�E��Nq�K��m�d(����P�b���滋�U -�9})�Ϯw��+w���z-��zQv���"0�U�]����*O�/���������9�Bb�^�h29���6׀^3&cD�tZ��?����NA.�%j=��&8�f�՞��̀8Fx8��n�$����o��{c��<e$Io���\+��-R_F��7���R��R��Ey�mR,��2�:]a�9^D��<T	~"��ƻ�Q���Vύ6��1������ڊ�S��z��e�]�N�D�usS�{�mz~����fҗ�-Q�d��7�-��&8�^��wB����$gI��5�[֧�&7��K��RnΑ�G���#�y���Ɂ8��D����Y�/z*���5� ����
�x�7�r��L���Z��r��"vXj�NЙ�Ij�*�'V0p�=7B��:������k�wg�����x�M=?�{���굆��H,Q��E/�F�W���@��N�SvjLGߥiʶ9���8���Z��(���c7��T�zU��gk�u�</�O�����&�(�k4���:i�IR��MM��xy����q#Jk�:����ɟRr㹁��*<Wb�b��@���M�j*��*~q���}�}��se�dY5��k銍<Q�םwr4���}��(�,��@ܓ�=�K�H9-`Ok��@T_������IUۦ�%����N�e��(���{��~{�_x b����p��f�P���F W�%��	�q�U' �UI/'��}�Y�ѓ�&���&qB�ii�����0`2
��% YDocc"ܭ���h�c=��6���#���å��4������W�Y�K����1"R� �M��֐��<���s��	.��?؟�:?4�����o�p%69�^yo3�4i���,�����s�m���e�Z�#<5Lv���^/�M����8TF�(��0�!�5WM�����aױ�D��D�׹���`�"4u���>:�v����oI=/�X'�J�D�h��]*�Ρ����g�	c�f�8����-�_�����G�o�-I_s(im`��y\��U�ə^q,�'�p�|{�n>�"
�(8~4��m��<�yd�sp�r��(�6A�ueb��!����U����Ў~��'	�!�T���a%3�����0a^u9��$ҥ�B�ܟ=� Mv�ȷR;�S?�� �JFC*N��6�B����:�-��9�#�	�X���5�()ť$McA��&�Z�b��|�K@��3{1}_^n�s�;��S8�$�/�ܙ��K����!i�>���1ڢ��Bt����&���x
hR �zˉ�����~_]�c�򽾠�ڼكݔ�]���G��4S���vs�����H�-3o��(5�H�c(*�'����8+�^x� ��O��~7�U��:�����n2�:�d��^��GM�=��>��3|g��_ܺ�bp����[s=�Xdr�t��zOZ�P֬�:�R֋����Q,����uW���������Q���#�]���h�T"���Q�_Yb����:��J�p{fQa��@�.����0�����@Y#��n���������y�N����o���kgM{����c]/Z=I�ydO4�R����/5��q 6�L�b���4r��A���t�J�Z]��3����o��f��v�����  �>U�ʆT��� ?�</����|��}s��2'G#_��x���|�ݚ�gd?�^��#Th�2��W[2�d���1��f�c�]hb^?��[M�� �����v��}��E'O�������ǩ'Iu������.�0/�6EL�팝��7���.7(dzY+��.�O����-טzrif*�o�ҍ�C��P��O@��}0��;Eй�w�.e�>���͵�1����>�7�:���ӗ?n?������9����.��D���c��,<���^����X�
J�˿��J�4c�Iг�+�$h,V����/+F#��5�j�%T/r^K���â��@��r���B��t1 4�,0dw��$�.VGؽW"�ksQ#���j���~��sn�_�Nd�4�f~$��r? ��O�m�#����=�b$�W��5<wٮc�I���Vq�R|� GƯ&5�X�X�;B�L�Š�w;W���P���G����0If���� =��n�D<�d����G�/����տ�:!�� 83�M�olx<w�֯�2Հ���y��=rt@��y�_�^u�H��Jm����a����زCR�Jț��z����J���~�ez��ΆH�k(���X�4P�;�/��:�͓	�*�;����Y�(Te��K}���Қ8
�@�8����ea�[`Re9$�D-�VLr�����+Z���Ѝ�?�Q/�b�%w��0�,�^mg.�J'g�O�0�a����e���ة��ϭ)pF��S�&&���T�Σ��sY3��1g��J��g���?Eu��B��3_���3�j�؅��54ׂ�P�t:���.n���E��t�6�;�c��G*��װ/��Yc �87���CM��Y"���}���Mu���<Sf΂��o�0Q�l�*��Ֆ��d�������%�ۀ�!���j\�=1�䗋��U��[�`�IfM��VVD�⡰xv"�v�8��zi���^�!mB��mtqj��W��r����/����%ޕAxZ���f:�p"���Xz�M8��Ld�xz2�:ņ�v��
"|{�3��q��|����(��d���2Q��Dh޸5ڿ�	=04�,�Rj��/�s�Y+MU3z����~=z�$���Ȑ|�<Q�j06%A���U�b�Nm�lS�t�(ea�����)2k�$�A�HM�ͫ�1�{�$��A�����t���� �0{��9�h^����e\��SG[;��9�2Z[��X}�"�,6���>9�Ͷ9<Ј�m��bYL���*��C+��;�>{�;�L�nikC[�+_K����M����U w��1��gQ@�`J�����:�����z�dMW��G.vq���,��COaX+�Gg���vt��b'R��rd? �ܺ�����S�w�s.�T�Ki�~�,���\g𖥲"Λ���	�'�Yֺpi����iBR˽
���
ə�c���_W�d3��&Hxy���"]�2R�@�G�4K��*���mM7����p�S���H��a�Q�����wh��kB���B;�]^E����Jc,�8Cy����PVi��F��?��O���jm˯XAd���{t}� ��E��{��m�u�/ ��K\6�uo}K��3(^m�FF��~&��@�K#g}G����F����;kQN�V�k�0F>�2����2M�x������q��g����?��R���fV<"�X`R�C�%��x�x�XQ�xN�c��hu�6�Z���}=	��6�צ��+��)��G��ɇ4(t��A�,�Q�q�8���Ԏ�6����g�7޴�NG�ƞx��������ăQ{$�L�y(�S�;Nc�r�e�+��ix��[:Ys����Q@��%�{b��DWeʴs�G����-�ϙ�͹MX)� ���x|=w��ʴ��'��;�q�B�9��v6�������I��1Z�������&��܀�Q�
��VS�H9�#�:8�*���H&ګxdRP��`�ĆJ���ܹuevE`MH^p����a�����ɇT�~J��c��6�4v��Z�"��d�n�[���E�<�3� �=7�zr��䵏IH�� K}��R����R� U!L'6i��'e�ʬ_Ub��HdbY�����[ϸ���J}_��vw4��r�@��^L��!L�]bV�y��;�[f�5�_C��OX)\�%K�Tg5��Ʃ5؀;�j�/;����Ǉ��\�5���l$��\��(�mY�}q��@���yf��k�9����Ԯ�[q�/H��g�	p�@;}o���I�'}��)1��>_�Uڄ)�$�W*�^)<�^��J�P�$d%'�������(Pȇ1��K��"�P�p�R�	P4	t��n��nT��O'f �H4��B��SF�z��G��Gm��T��Bd��pt�N'�C�8m��0� �;���zG�'��cJ��J���N'��H�`��S�\VX�o�C4�6E+��L�
?,7KdֆV�N�v^�b~	��'�iق�<�E4��~�%dVN�qx�[�b�i�[�Z�zY�n��[�X��#`��׭����-��p��O!��n/Q�_�P��u��&��(�;r�_��w�U-_V��f�n���X�^�8#���ݪ$�l�*�l�=�;S�U��C�SUWM+���)�z�L��_�cAK�ba�ڋ �^�	?��87}��h���w��f��G�"�:e{��zY=��un���kv����	�����9ˬ���؂��2����>!��A'�Ͱ���gѳ僻�Ľ��{ͤ|�[�Ξ P#M�$��{,?�af�G�F��:��+��3)p���,c�R�B��>&r\�)ׁK�J`)��7���]l��Q����h7��Ua��r�O���:-�Hn����:��e'�R�PH_: dP�QI%LU-�vTQQ���SCl�I��H
���(ۋB�;��=�2��v\:]�o�������^��Q��hX��@]/�S��ryl������8�>Q?� _��@����!c�ӳ���A	�������S�2߻��w�����>p��S���,T����p~��6y�;Tx�ԇ�[���c"��Ù[�w�PU0��N�(/½x���Hz��:io��$����&|���M`�|ec]Z�I��5�����L�ǚ�Wy`<LQ"�_8h%=ݪ��%�X�и�hsS�ƻϖd�F� 9U-�3xh�no>_�y�%� ͬ���(L�r���VH�L�����)���{5�.`�7xè��j���H��[>��~��n��u��D:��O9~ct#���yU��V;/�~�~�b����$õHi�;�&�	�H^9�n�v���Ean"�k7Dn�[�+���ơ#J?�鶥9{V t$�&�r���{�?_}��1��1�J�t?5�m�s<�ɍ� ��_�u?O��&�/�8f��9�O�P�G�|������[w-�>�M*S��D��T�7'������%'X͚��2�F/z��w~����m�|a�n���?�����>���,Dk�uJ5�qO*�gz߹�ѹ��W��#��ɇi,k�:��[D�Kj<�)OLEx�"�㤤F4��Bc��1�0[Q5��4L��e�^7���_����?mg�REbER>�w�bDz�Ė[�Wr�Z��C�$���>��J�+���٬?�oIq^��v:%�7?(#��lh���|PU�2,m�����c��T��G����Ѣ�C�akD�Y�p��ܾ��8af�hH&� �7c�u��$�޾��迗��z�j!�!��^�`����:�и�tC$�mY�d��CqT5�$�u1�_d%Y n�䝎IdN���&�ex�M߱�rk~��A�lŜ~Ts��&�GgFd=I�&E�'HBg�����(r�-�[���K̔�=���65��JR��;�k5yAϝ�=]�A$�f�X��rk�z`ͼ�R�I�ME�)~�l�<�I��d�.�LV��#3_D���Jy�&V�[�m|� �y�����C�����"F���C��;�N+u�Z��Q�H�ᄷ18
� =���hk�  �3X�^���f-LǷ��L��p�E+���H��l�p9>ǡ7|՛P�ȁ���ਢ�:���}
���o��WW4�.Jp���ߕe�i���xO�8	*�n�./k��jH�1lt�������D�CG%��Bn�C�ꅉ����/�=f:�<$]��Q�2;.�|.��] �i���z�de{A���X��4�E�}������y�T/H��p�P�I���4/��q�Iݭq�%m$T�GT��^)s��{�:����L���#Y�0��Y>�(�ON�<�ۺWU�ĥק	��90m+�]̚�}-}�=��������!����O:�V��k�鄼�&Ȍ�o!��Kl�4IF�0�,��y�+�ZȖ��Y]U�������!����o�.��g������.=��b�%-R�B����n����͡���*A �� ��@��Ѥ+\Ƕ��+q��M�RB�0Rl�W������n` ���'�?��mݪ�@�+m���i���P�bf������TQn�ͯ0��֯w����*Q�,h����_�}`|�ۼ�7�H��i�	���Q��wj��F&����g?g���2��]~�.�p����z8��y{Y�VEH���H�P�����s�Ǘ-��w�Ӭ���vV���`��d� ��.�Eby��n8jeZ�~JX�M�	��UU��QQ���N�i��C��!����*hWA����$S��ʲ���G�BJ:P#c�Xaj��[%2Ux\�Aɝ��l)8���bO�
4�� �DY/4O����=��I*���F��f�+�����Ī�#м�θ���]���*}���[+t�R^
��Q�(�a��b��o{ �璽��J�	��57��	�2݀�$M� �:��[=u%�����Ý!�����(j��9�6��X�R�/�D#CDǗOr�),Q�WnN����*|\�zK����qlڡ�Oş2d�S<]������B_��'��	�AM��?�� ,J�w�0�p�B�{3����|�jt��B-WG1�s��ys����K>!�!+ݒ�' QQ,���Z^�:�c*A5�g�����s�k;d��Þ��n�?9�����.L��2��ܱ!2�l��ǹ5�ҚX��.�S:fD���1`੮<����
EZ�_-�hF�j��Z�z���yO,�M�o�4�d@/<@��-:�磬��W�MA_�SӚ��מB��Gb��<���<���3��սj��r熫��L�d�y���ɬe2T=�W웲���ސO=F�����m�(u1?�i�U��:����	h{�YN�.R�lS�K�^��9�{[4�?�qHѦʔ��2�LYl��l2#���u��~�]��|����m;}�nyߘ��0��OQ�Gq׃{C�dmN��;HGW�]g�w������|�9��=5te��[�Ht66R�O⓶4��/��D�ۤM�����Q�5~�V��4 1�'t����57�R���_�fo*H�<��Kf2����h_ȇ�h@j��$	��j�*�r0�f��z�Ki��2��:ʍy��7��!j��nT�KpP�[��N)����tV4!�-+��l ?�e�M�Xl�;�ܣQ��K�f��#9��?��I�q���F[��7FB*���h��w�h�l|�gO5[��c9������WQ������n�?�iD!����u��'v��A�v�G܊�����S*ߎ�WիU@=�;*�)JJZ���'sς�"�z4'��G��:�^xz��7��D�n� "��t	/�!Q8SBCf���D�o�L<΁�m���=�\��.}5�\l{��n��J�Ʊ����ľ�㇍L@!V�S�:���bI���Lfx2M��)�"B�#�@i��# ���i"��PO�3 �0^0~���u���&��"����'��[���mu��?�x�u.�z�m�vE�N�K�_�<ƵL�uj+�Q~��#(��"������#?��p�8_�[^L挆�{HJ���J�p5��d�hri�{ͯ'���~�Z����S����4T�P*S�AIJ���?�;�,����4=fvԮ3�.�LS�����{�"�1Y,{�&m�M��N�j��1o~���U�Ӎw�k�Uag���l�0S ���)8�Q���o�>��!��v��UvZ��$��{�U���u{��{c�;�	�oά˫*��v�UU/�9�qP$͋HpZ*f���/��W�|�F?;��ZM��z������*]�K��Ft��5�U:'Hc{m~��O���T��e�^�}��c�2/�������֌�He�o��
k&�A�]yʔ��R4����Bd�:��Nm�U:O_ҙ`��E��7lE&�>�}�"�(�V �g璆��m����5g<�2
���>/]�B "���aE�#%xqq��>�U�t��(�92:7>�;3ه�`�)i��ﰬ'�T��^ż0쯯�Yw�d�U�r\�M����g���aqKdb{3ܪ�31��Zk���	��O�o������@Ҷ����æ��҃��T�m����#���?��c�Ne�������C9�:|09fG9�Cx��Ή�d�bL��x��ɘ��h��劒�������RN\Ö���M�5�B��ek�����f�E���h��ƻ���=T���&pQ�O���^��E`�ڒ�Dhb�6���;!�L��]㩟�;�:c�n�H�����rc-z�O����R5��X����d)�E���UY��!MT�~���~�����
�O�	62���%��T�[!���t�c�$�21�w-^nl�=�]-�y�`� 	ȩ�%��8L��s�����������q^9\�(�<l�]VH��ĝbc�7�����V�Z0ϙZf"�s����&�����������5���D"r�����@�˯�FO�Q;�%� ��|����\n�����`�{~�h�y�_	C-ĺ�D��掠�>���.�Q���3��4����!/��]N9ɡMB�]�����M��N����e���پfQty����� �]j@pk��k�ջj���%��)�m��{I�����	v��U���S%�޸��`�?��_��
�4ˉ5�	)���t.R�U��\l��zp�0��d�o7,������ ��[�u���/ ���u�-���X��o'w���^db������OЬg�G®L/�D��T��N���J�,-��4m��}�pYȭX+A�$pb��[S�t)i��]�UV�^?D�"�\��]}��*��ChV�Rh�M��eo����_��Omڐ��ꅈ�B%����:�<[oߝ�?GF(��X�U��9\���M�%.�.=$�3�����4Z�j�H^���}z��>i�����sJ7.
}\�gJTi&��V�
4�ڑ}�P��G'D�9��f���7#c����|�3a����0J�I����A����esO�"��H��g�Õ�<��OV�0>�3��5�����#țҚ}��(;�3^B[�Vsb`Io%a�Y`�.|��X�4��j,��5�h4t3<t��ݲJ�2��
._4��i6�ȴ"�?<oJ�|%��p��s�hzl8Hտ�9��o%��aRC/�'*�a��L{�I�~������8��o+����4��D��b�3��2�[����N_�̣�('����#kO��w$�Qi}���Pt�@�6
8�EN@��ۮ�2D��n�����2�EH��V�f�r��՛�D0O��1�5��0�W�1�ڌ﷨|Q��y���^����R[�L�o����t���a�=fVP}@CT��Q����}���n��h��y��$�	�b�Z�ٸ�p���k��3�j�=�%$�2�^�~�_�r��۝��8����i��A08���k'��M,c�����R�G�`�~�b����Źq��~,nO�?���)s�;Y���*�L=k�K��s0�bD:�d���g�-^|x拤?��)k�s�<3X[V�^��Z?[eչ+��fo#�pE���eb=���im�,j ����*�o��r�i���E-��>Sߘϼ��SZ�ƪd��9aVg�Mc��М�\�h��GvWg��.x���O��螚ޟFJ>r��4��o���'�۰}��r���!�͋p[�#�t��KIS+��=��8&�ٲa��ϻ)Bx��u&m�d�\�/u��=;!>��Ρ��iO�_��a	PW����9��G��/��/6���������~�9lM��B#�&o5�b�ϻ���j�,ɍ
`y�kub���f-g�x�JX��=6�7"�Ԋ�yk�/4��H�8��^t�ׂ?H�5������G��<�d���f-'������1�$7	�l��P�/ĎxܟRM���A_*�5��.'��Gջu����t���8a�	����q�C��4�x�"m�;�i���u39	�=S��2L*ʷ�E��j�WB�̱Ӌ�"�PI��o4����wG�IsqG��?Ma;����u�8~x�+�Q���*�/S�Ž���`�CcOʦ�ʍ����`Y	�Sm��ۘ�۟޺���WD:���1vJ�)�E�^ ݶ$�	w�������������j��ɟp���� �Q�v�Q�J؂8;����2#�
�s3�G"2Ű�`|x���F��kx9xe�����ޛ����#��r�{�K�Q9�}_D��Q�`Y<A��J��"�+Ê�;3���ts7�.gT�'�Ҏ�q>-����fW���䕻��ѷ����Rۅ��t����n7_r�~��>p~�>"�'^�rO��{���oB`�:*+�9v8�m�e�k0�gk�0�t
F��J�����!�v;�<ԩ��(e�؎���z5z�y��Hߤ���멩%�����	y==�N��e�a���c���31�0Ƴ]խT�A~d�f���KR\W�[�����-��lӂ��_^'aa `�-	��X�oW��ah2�R���`9������E���������We�_�O�^���M�x蝹���\SB�a��ހ���O���Gϣ�W���g	�������Y�N�W&@ϹZo'@�����s������#lr�|��fpB�� 0FZ�q�p���V��`d�'KX TI� �ztu]E�"�_D��է�|�[J#��!����<�c�f�=�W5<z}T�fK�j>��C"L�7^Ōʫ@�k�gN5����`�y�V�(�B+���
Ԍ���uT
�>�o�j��0�z`"�9>�OP��9��d��8�?&��!����(�HI�t��t���tJww��%� ݃tww73�0����~z�_��Y߷�����@g.0��z����@L^i��r1�p5�,�F�a(�[:
�E��U�´P�Ie3h����Ͷt��8yKbS34�w[7������S���R�j6�ay�^[�����ۄ�:��2J?(�$b��������t����em�й����8sm/l��Kf�l�\[�1���0x+��������.ئN�+�b����jO#"3�$���e��[}gU�4@Wi��Cx��)R#�W�
h?��I8E��xJH��Ă�X>�;������!3��?bX,w�Z�.-y���������!�[LW������i8�A�	��C���;-��B�n�#���X��&]�f��|�*G����9�Qi`!C���C��|���ROϕ�L��c_�7�?�>��}�PR�{,g���z�}^�F��X��x­�qn��^.5��)��ӽ�Ī
��$��eI4.�[E��a�	�rA���
{�D6��E�p���������.�iH������ޗ{ |��s�C�b��P�v�9 M錅w�3��;�x�T�ti�r�\tj�*����j	�����h/(G�D,�Gi����R�v`�XrZ�Z��˚˃�z�\�{-��-v����$����>�֞/a���C�M��/���ærl�8n�}�08oM^b�ꝥ�ּ'�#���d�R�'���}%���؏%`To��LƋ/�w�Q��&��4󶣯v��0����ks��Y�o�&��*~��,h���� ����$��lg�*�)�{RD��mU�S���r�ޛ,a�R����??�w�Z��)�GPy���$��-3��lV���X���w?�%M�bi�7�Sl|/�-��X�����	��K�2�B�,�꺆���vzl�p)`	mD�r��nG�L,r�?��g�y�Q_��N���R\w�EVP@�Wm��"� ��Xߦ�)��Qg��/�o.*|�z����6��g�'^�\��_��8G��\n���O	A��Y�E�ȯb���l0��R޻��R*4��22|t�s��Aq{�&1/L$r�:i��g����L��]�j�cYjU1�A�0��7L�(���!K�s�l&��f�sY�t(\'g�M�B4�_�"�6]Up7»��&��\�s��e�lK3����S�N*�R)m��Q����ǧ���B߫�ʵH5��������ܾK=DJ
�O��`b��͌:}Q<��zm ������ߴ���`z����ۏ���8�:y�'�H���N5��G�'{9�Tg@亀��3��R�����hD�37/]��N��MM�/����S�.��*��X/t�#~ɣ���3����y����0oEO�[fx=�C	�ޓ/����"g9��M)���7)G��*���>,���"`8������<ym��I�������e=�����eF0v�ҙѻ��wt�Z]�Q��=$#v��s����`\�r��ۿ"LOz��s;;�ޭ٬_.�� �HW�E4�zE k��m1��4��!8U���7����J�����Ao煗;
�nv'�<�tJՕ�$�0C�ԃ�;��^y��w��Xi[�2]�!ю�/ƭɍ7�C��x����̸��B)0����z%}h�:T!z�m�L�ƒ��g�/�����u� %_��0�K���[Gыw�4:���0WN����G����h�j��k:��7Mn������ee=���ֵ򪭟��v:]�{P�P�Y�gi(�w���v-Ckr�3h�{���}��^w�n�9�����SRTY/��/rCq�J�mE��Q"?;Q<L�d���$��GzUۛq�r�Jۤw,��K{ד3sF�G!��x�E��øuu�B����gvo�u�f�"���Ӳ
п�>{vETt��*"%�դ�;��0��M���t�a�D�<�_�Sr��zGoڃ��ЋF9���Ani�����q5�,qQ��m���igV�h׭��[�/6O߇��.G-� �=�8c�;i�U"B{���R�1mq�r1wнIp<��8��z��̇MhD�$�E{��M�T=�$n�r�K}����mI2u�DM��;��n�����ĉ��1�BY0�\{Ǉ�:���^7'���hG۷��3��~۰�X����M�(���<_�d�ό��V�ilK�W��	�a�z�<ob;�_䂟P#H�s�`��m��j�u�v]�K:R�qj�E}�.�D��U>b�QG�&�xI��4�c���Z���|!�Ȭm�ٳ��$�lA3.�̎��ig]�3kGܾ2F`vO�Bi�Ϸ�K�H�墡e���i��I<���'^���O�.sr�sJ�"�#s;��g�%3��g���5~�8x�@7ý���3�Ł��=mi�T���i��7����V��OT�A�fږ�L�������K�D��䎩�e�$��Gp�AtcT}�(���c�Ÿ���җ�ѯ��ufSh�&=�Y�aOx.q:ɘ�.�m�˿��v]("�Hs�Kh��&���q��[��ۇm|h�t[�pn9j/V8�7U7�>~螵8����������I�y���WX�L����7�3�k��g��B�>_��)��YU���W���W.�y��4낼.��l����
�����vQH����<,ꌿˉ����Y�y������"��w�e��ٶ�x<����F�_M �јh�g����xKN����^J�ӥ��u"=�\�[ �8B�þU�[+|������x����:�b!����d�Lo)r���N��*	�km��B�G,��sU$�쒐~��]IB��[72}�E��Hp�}��+�c`agpv��H姭�0�a���Q��������-��ӧ�Z��%�M~�.���������؄W�.���m_;+�/keWV�Z1_��y}c������	�c߳=�Pv����-���l/Hβn�o9)<yRB��M̧?�@,��������x���R�4���==�4�=���ys,�����Ĭ���1�A���k,��wr�(G4͟jjۛ�J.>��jX�On��o 	ew)�2�l�����(] H*H1tk�}�*����.�2Z6�ğ74� f���������ط�w���3Uo�!lS�8r��	�T5��w������w��lI����k)Q����KB�3�0����U�º`��q�z>E�夷o=��@���F�9k�Ϣ��]X65���J�~�$�-�3~n4����b����XY>���֩�O��@����d�6=s�;Y�8ߓ�q��|%�	��H~��C#WȮ"'̆ZY��1�x}��,�I�=b�P��^Y��$z�O
��ү1냪�et�����fD��������P5����<�S�~���V����0�}N�S���~�$�_UQ�P�MXl�0��&?/D��7���'�E��L��jyQw�~��]�޳�&<8����r�fG�<�P�9ц9�GgOj�}&����L�8����V�%�Dg�%��/��̹!7��H	��+W'j�9��吠�RO�省/�o/C��_��9����v���9:���\��[��l�nx���f�Km�Ұ��θ�J�윽�Zps6���~�0�z/.mX���B-��P��K8��w�����J����{�@"�e��k�D���'±��۵�V�<c?�W���t����-?��|a/'f0�)��>�F3SxAf'����4zzC#�U~�r���������&��[��d��\bnU��:�N�0y�Z'ᘓ�?�M��|�|�a��È7ݧɞi*:����>odE0������y:�~��L=a��<�a��4 eC(;:O�k-
�_��L?�Z��[X���W���j1��ʝ�|�]͡Q��h�
�߂p���` ������/�J��!��C��u�������9&����kJ�>�s��X��:��+��T�-�3W�&�0���7ǥ�K-`��7���R�y�����|j����f�V݁��'���;]��͐����
w�� �#��������GWh�m"�u$xŜ �<(��>ҎGM���\����]#*�vQ>���J%ƌ�r�Q��d�^	U��� ����H�un�{�^�$��yE���gE�o�m�7A~^˶ߵ"�;����ON���%M��_��\=T	=�R(�i��x�����N���f���,����IX}�@�s���y�"�͑��X���vS�h�q�}}�ɼi2�}$�#��y7� �}8���������6��5�o6����+b�RF%�7�GE�uَ̅�?b=�:8Ē4B)`�[`�z�������-�3[(�*V��z���b�������ͦr#�!<�����L�<�`�K_���f�V7̙۬Gg��/s�o2��TȲ��-P���_�&^u����=��P�!��Q��D���Ʃ��K�N7��0N`���k���E���숉����Pr���w����.5����Ұ2�:�#��ʳ_d0�1-�����ph�S,^�ԉ�s�M���"R]B���3t�e��<��V�Z��U���R�cmj�Y=~<5b��B�xl81�N	��G	8d[>}N�ݮ;���6f?ա\.e�~��&N6�&v���54��%�j���,{_ɿE8�b_q>�pb�8Bh�k�j������u��F�d����P��������/K嚱aJq��3]�m��݆�=�bu�6oyn~I�Yt�J1g��pr#͏�)]b�3w��Q��X����0C,�^H3�gN.��ؓ�6s@��J�h�<��OO�=
��)�v��B֏���ּ������X��-��z��}͓p\(�g]E�;��$��L�u�|3��P��穲�SR���i��C�K $�׼�3��h���u$�E�s1�{�����q��0�dF�Z���1��Ѝ��5�Cǻᦒ�ض��ű�/�-!^���M�S4Ţ	I�H|�ƛ5{O��C5W��yg6R!M���]k�%B�N����)z/{����C�w��)�*m�Yc��w�g��hv�io�����A��g1�����$�o��
�5��=��-��Z��!�|���7}������-µ��M,����lG�n2�r�.����S)GxW����g8�B�Au�:w&N*C�=j�3�Ju�;�uZTx���4��%���t�M��4}��xÞ�ܷ�( ��M �����%�ݖ�~Y���|�+�)�ꓫ7�Q��G�a�Iy��5�����5���}+eR�x3��Y>R�D�p?�M-�^��YNUO���z6�%+��''#6�[�WW>�4�4Y�,Y�e�)sYC��3�ظ�K��i��X/�Ev�f��c@�P�������O�{Ϸ���'�Y�4����qsd~N6Oܘ�|ˣ]@�{U���\����e�]*��745�?���K��n�.�ѡ�|"��������rH�I
��?�z���	��O�Tv��Kx��hO���0���nI�,�Sj~���m��bd�'{�sx��i����5���0�9e�3d��L�%,�>ug�Ӥ��β	�<��@h����^���$<d�{!H﫭Vq�����ل��Ek���}N�"/#����{�Λ��P�7�F�X��_��&�QV2�������'�z�܃x/=�{�#�7d��x�gaΉ��7+j�C4љ��|��~[�u�a����F	#9~�4���ul�{Yguf���#l3q�X�x����K؋�5��id����#/u�H(⟯�V��7RW�$q>m��
|��`�E�c5�W����ջ�6�}��`�����z�W�=>k�1���p.H�R��y>3�IO�VՋ#!�s0=ش�j�}Ӻϖ���r[��&�z���[�Z�+���k���v2��왳o�l�� \Wi{��i�y��D\7�:G���'��d�:Ud�|"�	���SQ�ýoӬطx5�%aZ�M��q�I*c�?��!�e}ڹnHӱ��n�פ Hp�N����v;Z�]+2����Q�Z� Ȟ*�x)��`λ���)j,�q�hj���Id%q�-���_5��\�'���^�(Sԕ�?��^Z�m�Zq��_A=8Z3�J�����kH���[ʥ�~�yF�j�o	"���N1����r}F��;��-S�Q��d^>yu3�	io��[x���9h��������r1�s�z��eMOO���Y�VI�aj�b�!�6�jkJ��@��'0y��H��3zZz�|2pM������$}�k��~OPh�u9K��J!���˘�ߦ�B?~\�b l�YEJ�N���|xo�W����"\����82U�[�[*2�Q�΃^�F5A�Y�U䠵�"��~_g���������S����Kt^�ٗ�N��d�w�#?+����@}�����8:4�h�ѕ �������o"H�$�h����.,��5;���,֒�q#�����>��E�멑}�$��������gg�_���ࢄo9��ަIsp�\��]�[��UT�qx�KAb*
�8>F| ���:�4�l�J�}Y�TgB|��8j�����Zu~�r:��s-0۾\K��������ۜ�㫫m.N�C�!�Z$�����~�}*�{j�෍��|ͳ��V��9;l� *GMW�y��=H"_UC50�tl%nK���{0{�^��sOƼʥet�nɕLr4p�?�: �c5��+�Aۜ d��*˓vh��VNI.n`�jae�����5�Xc��.�nO�c�">D�G=���e�\�i�>����������a�\�g��Gk��Ⱄ�}EA*��p[Q�=]u#�.j˧+���5�2�\�@F�F��՜M{���v��"_;�K���$���n�N ˎUQ��!�l����Se�����D�����P� �!����ye/n��S诣��7cK�a���#c�- I�_��{�ر�cnf���VCI�]��F����K������tB�;��[�/=�H��VW.��ܫR_�yxu� �V[�]X���5��_�>��'�MU�??G�nd�-����~�8d{R�_�����S1���:cph	�W�G2���Ԭ��A��g;Tѫz|��l����Ys�I�O��|������?"+�j�}����-\�5����{�����s�n���A�%��VT���-J;��F�A|;Q�,x�X��|7%�8h����^[G�LZΞ�p�EZ��Ȉ�<�H &)9z/�{����f� �#+�'%ʃ}l3����}�JK ������(-�tOi}哏�Q��+�ő9�@>ވ)Uś9�ĿW���`�����<� `�Xgi��x��?Wn6�X��3&�}zN�+xr	��^�׵(�sσ{\t鉳ʞV��hkz;�)��d�.-&��:�N|�*�>�K�=B2��lj���N�uTֶ֙@�+���|﷢�c�O&����Ȼt�F㑑����SZ��/tVY�~8_�BSj��Ν�5�w�L��J�G�;�u۴<��3���:ϳ��֮x�z����>�OzQ��=U�����1�����F[�N���{�?	�|ׅ�J�"��(cϚ�I�&?���xᡠ[ue�x��������$��:���C���b+s`��R8T��u���"�*��n��@�T�ˀ�+mgֶ?�xp̥�j"3Ŗ��+��w�b�ˍ>�Kce�V��,&�f���C�l)lx�V٫���l'!7B�����5��	Y�F��"b��K}/"&0�|b�`:�KVj��"(��J�]��k[��D(�R�$���'����I+�P��߳��Y���`�M�P/�l��H�2����y��)�����Kz���B��:�6�L mݵ6��2m~}��oJ��0y޿�+����r4!M,�`�u�q�XB�V.��u�e�u�l>+��z~�\B�����qMc�3{���h��E�����
��p���'f9�ʅw���q�A4���-x��^n;�,�y{��@aQ�#�h[�%�O�pn�iP�T�և����x�����sF�������'�W]݊�^�z]�J	b�&xE� Ѧgʳ��[�8���5��4Z��$�G��ק�99����Z7����}@ΐ�)%"�Sa�+��>��N��0�d���0�(���s��CϬ4��e�B�����4�+�$M'u9�x%~�R�i>�=�U~,��鋐��Yn������,CN�����{I�rX
�y�&^�X���~Bo����FPl�D)������}cm�sS���t|GS�����p��M};&�����R��s����I�#��)���qn���s� .쉤�v��4$^T�����+�Z�^z�0 w�j:5�gk�sd��<��{�!l�(E�m�p�Hv����Y_�l����Snjog^�^<�z�c���%��D�\f~��"�@�ֆZ���P(�_a!����9�U9'��&��${FFU 8��\7]ז�p�t¡*=���1Zg��ko��jK�s�\�u�Poz!ۢ�ǍO�c_�z�5���n�	z�*~���,G�֎H}�>ť�3b|��{'�M/�xo`������f9xRe��N�����qt�+�b�*7*�2�$}�T$�b�k�	 ��=�YE���e���[Y�e���+}3�=��'�8�ٌ�ѧ��E��>�9������X{[�d�5����z���U���'���T'魟W�4l�ږ�dZ,�\	X*I��Aj�����3�G*ޟ�NXXT�_��*&
���X�ca�P/��(�}m��ڥKS�5�>�jY�م�f%bo���ܽQ����+ 7��i�hM?x�V$�`r��Cq|�p���h���Q�m*�����]A8�����Q�dz,p�n��k���@�#ă6}�_i����ZXKGxgF$'�mɠ(Ϸ�Z�2��A�f���]�{!u*"͙�`
�*��G+�������ic���WW"�G�o�L�L�|؆��M924��TKY���3�����(���+�a�\S�r��Xhi� }���a����<��*������;�Ǯ�b����?<E���f���z:7њ�߿e�ƍ�<@��O47�r�A	�"�>ș�`�����Q%Q�u��֍'Pj0-�4�]�m�iC�����r���'�J�!m�,ȁ=1trM�ʯ��K���xop�TR�x.#�m�Z͘	���vn��gY�}����zw���} ��z�\i�f�QU����0�b�\��w�5�1�����O�]��0�kA<s�&i��щ+��P>��#�s��#�m�Pdr�;�.�-��5k_>K=ܩ��f�p�ds�z���A<!5��_�?E�(�,�4_�:)���LE��8�6^v�P�Hh���H-KR'q��%����ha�&�pOj����rf˱Y�hr6�줿�7��}��R���J!6Ŋ_�_�?�qGO�S����� ]'z��X-��	�Y�<ċ�#��p\�a�o6���)�m��e��K�Z3{"�}RB����Đ3
�seH�fe��gY��կ�E������5��0=�bX��I��@/�����,��!�����C�5Z+6�4}8�� 	�{�������N��䁑&�z�I�"�K5#�eS*1��d7��z�2.��8���\��/Hb��3h��f�"��d��{�Q��=�ũy��&T�vx3Ǒ�]_�`�����;h �g_
�
I���cU��rª�oZ_��0��yŢu�&vm�k ��n�]q ���a@?Q.\s���Y�W�+���+��{_�w��:&��x�-:nEs�"����f!OI�����ʆ�S���zRd��R�������+�Ʃ��Ɔ��׼�[/7�rg}�'�(�f�n����(C�4�,��Ϣ=1߆�V�Vt�-�΂�u�Qi��V�T(��w*��ͯ���@K�����Bx��sv�t'����aN�ݤG3f=��bv^�!>}��[*����o3��Yd�(�K��WS�睷'��`����
!��r/N^��s�DU��!� �1�����u�sJ}�����'_o2*r�ͺS,\
�j��f%wGQ���3�'(F8Xd����&M��M�AK��}(�ᛩ����]��z�ɺ$s~�k_H+���ly'�#3\�r�*y�.�:�T�ԕf��+T�㉅�瑘��h��c�m�24s\4�<~s�5F��T��S��`Jl%�2ZI���gR��x�����x����Nmu=3����0���~<�X#���,ph��XX5�T%�m��f!̚����C�}f������
����~qOe��zdݒW?�|�N���s��;SUe�r���D�ٛ)���;Ko)�h9�e�DD��0��lޖ����2�mQ��1~�'�s��[}�Ň�����pm��>��+sWCp�w�'b)�#TQ%��w���DM~⯂r�8�X���6���ơ��D�J��w�>�H��� wI�����ϟ����R���Y�ܮ=��L>p���:���xGWdudT�dl�E����u�itHBb�qX?��<�GRs��Sv��	����9�Yx7F{�G�F�9X��3=rH�zk$���;�����\X ��k�jܴB�f��ɶ�X|�#�w��p�'�p�y�G�.�GC�9X�u3��_Ge��Wk	�lֳ"�=T���c�2�)s#[�ݎ,�z�ξH��e�V�4�2��#�"��$���_�Ԙ�@��U�!�j�8I�p;хi��7v`����&����n�-��[���7g'$6���!o�Z�D�M?�$�y�<}ivI�+:#�[kklÄ#v�g���[M�1?����s�y�{�����hWt
�
��Y<�v7�r�������.���-	�,Gmnjs����|�6`>DHUhJ�5��&@����[T��0�8(�W�Y7����g	�IR!Hv�.m��]�;s)�W�6�.��g�\[dD�D,w���b�N!�,oPe�V�j�'�\m�;�l^�=��������^�޸t��!��Ɠi�~�g]�M*$�x3��Ñ1X~A�LPF�kO^^~|5CO�B�AFv��G첦qTL��
�>���:��U;�T�e��
 ���'�DA�s�7媪�.<��	]�4\N��m쭒��82
ګ^OW����S
��,0%M~HHd��x��[K�,����S�1�Vy�̌��-����Uw��E`S��|m��U��S�J�Tn�d��7>b�Ga1���5��/��Zt�û���m��]�M\$�Z٨o�<�LK�;������T�cR�嘊�z�����]�L(��!UW�l���(-��?`��4�=ۜ|yuumQB^pi �v
��j�Δ�\Ս�3)\>4��^��������v�����,������t��hQ��N(�OG�#e3�r���z"�D��� ��J�q�n����h�x� �pl�z���i5�vZ�qt?uHEO��U�].�-�LZ�U�숄%/�K���D�]�����JmN���I�:��E���6��,��/�w���M3 �F|�ytT氄~IV*hX�\HJ��u�N�̃i���}�]��T����y�Z��?����9w�D���Ќ���w̌�@'/O��\�7e��ŀ��V�$S.JU4W��S  ���'/���Q(���)#�j��3d#l��%��1�tu9�j5X��ȍV�o��8��y�.��A47Hh��J&#�"Q9�!^Yf��MV�$��oj	�]�3|��>���C�0����Y�.�D8p�n���}���Nq���;?~0�!�H��2�[���ǧ��\`Sr��U�������̏q����zerR�.-+�8sZ�2^�i�����X )~��>n�<���]�=[O�
1?�H�ԍW���L��,DM5M�ǒ�.%���]�%�:�o�_|��۱�ɚ[^nk�W�U~	�G$��^�2���q���(�5Dg��t	s��l��ӎ�&s��1�?����965κw���̨��yY�e)$�=t���_z�
��P&\9J$X)W �K�]Dƅ���`��)���������|�a��=�;�kRwiKi"�om���$F�&z�ݩ�Nic ��Z����'�E
E)l�S��Pr�e�Q����?#�S����2�~�o�9"�G;u��Z�/h��azB%aEe?V�k�m�I�̳ȁ9ú9U�E�K�a�rh?�b Y��F/>����U}����]dH�=ҮU����&��7���	O�6\� 4����^w�1���J-x�fp�4����/3�(2j�o�݊C���4DFh�� TI+����K�]9J*Y�3�qw9���ƫ�2M�B���o5Zu��8�Ց���<7U�Qo�h�Ñ��d[@�r�*�[R�5��*���ȼ�O������E[�r���`!�䋫Cv92�]�YK7a�:��
����~�������{�BJ ŰU0DB�]���t��h��b�����+փ��!�?�?�bR����u,���K�v����0��#˲8J����V��e���@>�����F�^�|����:F�r���~�S������͌㨇�ڧl���V
�mV{H���M�5�,�tpq�:�74�t�s>�|�b�P�Jk��y]/&�?�������9h�J���O����������W?���n�/�~�ܘ��T9�厊w&3�=�n�(;/+k�V��(�<��.G��]%.>Ĕ�
;Sp�mw�/���sV�r�ӗ�(��tM�'��Ya�9�b�#!!�]�o��Wc>���,3�YOJí�����*X��Φ|���sm��͈�}���ы髄��/�
Ķ�b��"�m�������
���n���oӡ�y�=-��F�"�g�����/d���%6�����(�z���hU�Yr���K�\�,]v5I�܅%/�+�~���0Լ�8L�|���}�E���F}C���s������y�-֗���9�$��<͂5�<�/X���+-��t��߱u[��z�ͅ����_6f�����w�5>�m��r�����X^��i7˥qc��r3���81l{w�.B������w����8B���/�qց��\k�d�'�k2����*--��^���bv�Ȗ�KM�F���������p�}PU��m�Zcl8�Ѐ��Hl�d2~e�"��$z���[�J��/��buL�{{�p%Y%(0�O��5-��}�?$����8��u�<M
��_$��T=u�×}�I�@pNؔ�_N�#b[�d�i��3q���4�O�=1�+�f�#��N���x ����~�I����ܟώQ�E�4��u�����?���<j�䘧B�2�!BB\Ы����9�-$�6z"�f1�����g�,�ym�'�t�bVC$M�=��
J5|��5��K8��X8�wm���7���1=�<kv����9G4� 1�W��м�f��ȳx��9P��^�^Q�"qk;�\�{���)�r��E�eԌ�]޸��3#���S.ӱ�(U{��S��-4��)�C|]
k&|S���ˍ}��lo�h�$�^�Nm삘GXx(�E-���.�Г?S�,7Qn+�A��r����ȴ43�#g���a�(%��!SO}�����x+}��xx��&AC���l�PPe��}h(�y��UX����F9+$��a�h���U��`����
7��NT@��)��r����Xж��'���'k�s.�)7��^-����������3�+{���dB�����Q����"���H�h��8m�{����\������ɕ�+mc1��;��mng%�g2�}:��8�'L�[��Sa��B���R'�W*Ů�J���|o�4�PX'�����.|k*,)Qӯ	���)�15���I�jdr&ڌiW�6:u��%.,ݭN�W曨获y��f���ĕ+9R���[���q�C�4�
�'�+�(�7hƆx�n�:'�$����׌�F�m"4��C��;�{�Y�n���-���ϋg�Kn���۪X�fQ��԰������f���f�ӷ�)���{*u��鲰.�h��kk|�5���"]�F�Y�^�y>�-˥mzM�F��� ��_�g{�1�&'1��旾sA��7�N�"ɀ�o��iz/L\���M�y�Go.u��ʻ#%�G���Z��z�*}�vp��&~xe�.�b~��;m�M�C3�x�C-�Pu۝�W�"��'\S\�z��&F/�nՓ�x�TYN�jG64롦s/Bf��iB�����q��Ƕ�� `���Y�x��z�2#�{<��qNzt�2��c�`T��s���g�>m½B�Mf�+�꣊O�h��.۝��v��!I�%־&��7��e,�\���V�������p?�N[��$��\�"���v��h4�~�`�q��=����N�P�Y��/!�v�5٣���z�ez}��M�(��-^��my�]�wc��[!ޚ$�{S��<�o���/	��/���3���1 ��C��[�a$G�#��knw�r&�7��)j*�q������Ť�� '�����}55Cf5̳/7bZ�9��Ě��U/J9 ;��B� ���� ��Cz˳�_��5�N����+)[dYC7-�nnc�:wv�;Dnb�k:i#ШM�Yl��| 3��4/)V��)�5!��|�KV
�Ȳ����������pR��r"����Z��C!�΄�(З�͢���7?��F���z���Ug(71ǜ�&�r0b��i��:rYGC�W�ɻ��O<��?�[[ !��j��D�y"�BS���+]���ZE/�L�DK������|]���O^LO�t�'�q�^�l&S�-��sV�X)X�f���pu���k&U����=�o׃>*"���/W�c��8֖����"��� 1vl��z.w���W��G���pF�T;�t�\+�H*u�������[���l�3rP5 89���bm��� Xp�[���Y;�gKlr��M�r	��d��W]���3ͧ�����[Y�mn^�Uί��`�+/n!~d�'X(�O1�Su����T`fP��x�<�4N����mA/VW�h�x�&�Bb��3�~�N6�jB��ƌno��6[��E��\�!���/ɝe_���h,�ƈI��x��i�߈�b�mHh��DYPP��K������sK��чľ�P������A�P҅��rV!��K�ioNG=5�gs�Qhh���'㬒�ͳb���m_�(����J��i�%*͔F�f	i����"wr����Y���ڎ��ԡL��m���e|hH�񶶾���[�b���0��Uv/�d��ΗW� �����+:��n���=��};�N��YG˧D�����S�b�Uϳ����'��B+�����7��{p�,:W0��7�������9��T��6�y�2ֵ�b4g��G| EG�M\�\G�������/�!U�h&�cMy����#S���;�|Q�҈�iv���&�&_K��{'��d$�}:��}Ǡ_N��8��GS6�c��ʑ4�%�EӠ(iM|��kX}��yM�r�4�qVF����[�Az�}'jy
��4%C��AY�,��O�o����O�v˧+�z�	�J�����u8
Aed���a���1 �+��᥇��M�ށ�c��/��R�m��!-��b��uN�lc;k�7#����8i�e�m�JA�����h\�oӴڦ�P���-?K	5I�d�f���@���-���@�t�qnw�G%�|գד������-ݧ�����
�%0]�+[%1�����εv��n|�ގ��U�^�U �	B;3eR7:*?g>�}�u�<��˺�����	ā_�J�U����k�$�4l��6ն6gԴ���1+�y������ǂ�=y��k�\G �pǆ�f�˼ſZ����n�g��x#ȟcW��x���p�p��ɇz\r�N��K�;�F�y| y���4����TVH�TW�8�؂�,��f�ț�>X�,���������r"��[�S��	���%.m���%/ϧ��K�pj&�#_Xu��u�â�"�R�}-�Y QX(Mݿ�تm�����`CQç����p�"s�9<������Ib�jޓ^��IsIڬ�,J���6�K���M5�c�ω���3�_"���d`s��&��/�ʟx��E'��<�5WZ�s|�>a�ʮt���]���k�,����I+���VP�4B:����1R���XJ��r�.,�b�x�
�5�˖��6ꂌ��.�G��q�<�?5�H�Ev8`d�+-�B�<��H��8`v��|e*�s,Q�p��1�3=��!���}vz(.���`���$;�Lx�hL	I~MbH[����+��^߰==%)(J
H�Q	i�fJ���c����ь��3`�FH��QcCb0���>�{�����~�羯�z���VW7�:rU�+x��:��b�b�Ɖ��5{!vP�'K��Q>.�e����%�Ek�S�A�ÊW%�_�CLT
t�_��E턡M�o����	��F���Uw_�&�|m����6����4��ܠ�us���v��5P8��{X��?L ��&0�uxԚO�U�C�nY�Q~X�����~[�V����/��;o����=wpT� :k;7���6} A� �*4��[����D9)(��La����7i�B�n@q����\��0>�"���Q�j��Tg�_q,���;ͪ)F�r�Eٌ�>��p����m�E�P�kT�E;�v���6tY%�N��N��GǮ����ue�,OZT�%U��x���=!ϧ�x'2���^�?>Q������	�b�(j:J��a���@zلW1�U�SX����N������]��i׽�Zvz.$��rJ�e�i�� �l*�1޻=I�R?Ϋ'ζ���R� EQ�Y���� Y}PS��bd�NNN-zq����-)q?�r�G�?��\A ���!O����)&z�].�z�_?�H�%
*�=r��>�"U��}���u7"ɗ��� ���na=E8����<I3��ǲ"j��0z���N�q�?���-|��/��(UuO�I� ә����C��`��P��$G�ʕ�~^L���?�_��Ljd���S���aa�C}��ʠ f����vv������	�=�?�S��d���,C��O�� ��xaX^zV�R>"��7���efT	��RL����o��?��}��o
Z��u<������L��6�Q������o+2�Sf�cSW��ӎ6�3Sk+�>��a�[�2�͔��v�y�S�!�����c	���p�����`�WCeq[������a^ �j��8Y�9"��#��s�=�(m�C�*��;/V���1�>Y��it����RN+�E溻2a��h�S�5���׳w�D���gZn���ތ���L�i%������'ps�{1�<�� �ء�il�B�8�"ۃ�z�������c��ΐ�Q��|MB&�u�}����r�dm���v="�U]���,C�g�R�����qs�G?�ɒ*�^P'�x	t'S������'д;|��{U��?��z����F����{���$��I��V�Y+�Q�:�������O)%�\�n��[�.�@�v����i���8ό���ƾ	�{���騵u�C1hO�ԋ��c�(����TFZBC�5�'zϭ(�[A�xP����|?�Q ��畟�sr���_�y?#g˗F��L\���V"����y���[z�E��=-��d�!�e����� ��PLo"3�e��>/zǀ�Á-ŗ=V���6�Y�#�נ���!��m�S�S���9@�Am�Y������|W�C�yײ�.������|
�YNx ��s���l1���J����J�Z,n��U
�gG�t��f�O-촕��J�I%g�����
����d�1gnJ�g��ۉR�F�9>�E�����U_NY��%k�2�:�%}�H��43�Q� �}���s��i`�c�W�dP!�-s%�sP�}vbK�ה�(��� R33�a�k��pHz������G�O��M8�-Kɞ:����pD�oK�]->�,��� ¾@�5��y(���/1�����.���K�d�Tغ�6�>`�
�sy����cC�����#|%t_���I��Q���ƾܘ0�W��M�
<G�w]����
�_����i�Hx��G���hQD�62*�ef�\k��{ވ��q %�R;ٛ���H�Nv��1��KQ�� v
W��_Y��;#���+G��+��9M�Y'8�x0�H�@B�[��+舃;c��l�[��(x��޻��NѨ��޷2c�����[���g����H~�rhu���w> ���rM��O�����g[����@�z�x�A{���N���kC�FS2(�0FD����ߚ�ۅm9b��+�����RyQݓ	���ó/�*9�ꐌY;W�`�������ڪ�J�$�Ҏ��pt�2hJgWQNP�"�n3}��?[����=z�����M��%ԁ�x�ֻ��r�����!G�����5��E~�^B�8_���0'������ྪ��>�������I6����Ш��0�������Q	&�?��'bCF�a.I�.����"����>��|>�6�2�{�����4���X�M�*JȂ��0��U���^S��VU�2Oe�cA�u_��i
q;r�����3%��<U\��ܼD�R9?p���2��'��\�����W��4��%b�zG�B�a��Fpgnj�����[�JF~�����H�U[]��������t�	�c��[���G�!��`c��t�pi�Olu.�	�|#��%����P����pL=k�T=��$�(茴=)D��\��;
��S��z��z���3%"��9��,似]-��.��ZP]�}IT�ճ�#��4�/�q��k9s���#�9�B��A]������Y��B��GJ��Y��)�๎�c�smbn�Kx����,j�0(b>�ڼ�x��z-mՠ�_&������n��;����M�DQj�g�5��$��h~5�����U���w�YZ�?��1,;��u�Ik6{��5~�Q����+%�eW�:�y'�6��v3�`O�V�6oz��@W���?������p�ކ�T��1�I}�c�_9�Vg,�=V���K�L��oA��lk{�c��F��e����L���q�Q������;�'$��7 _d��T~�@8>p��\��R��ދ�	YvM��Ə��C���&	�@|v�s7z	rneB��9J��#��>`�z��w㴐tg��c�Vu���$�[t��Ϝz���f��MW9�:�	�R4�涱�Э�"̲چ	w��Ӱ]��y����)��^��zX�(Fg�`7�EN�����әl�)�4qL����k�J�s�I��,oQKM����/��f�y��:h�~�y"��l����쟩�v�Q���%��{c]7�o9We��Gu�	�������#�'�+��O7��$
����T����m��6P�Sn)�e�t\Y���a�R��<�O�}f����u1w�}1��J�%�'ٵP��AqԘ�����A�z���`)`R��$�j=eS�ytm��t��7\#�g����y�YfӬ2���9h�5���I�gU0c��tvb��)���$�T|����wu�ؓ��;��L&�%��乃̢i!�R��!��?�)F��8�6j^���M�Telp����ie"����\�c�y��q����D+P��7�����/Wp������ͣ8	I�=�� ����ke�*�~?������	��쳺:��o�����7H�RJ�)� ���/���8�Ɖ��kg�[$Zl��LI�ȧ�>D �d%ʗ��6��:~ N�=�'�o�<X�R;�N��;־�'-�b�A������O����4)��Y��E�w;w�u������߇��q�N��x2>������(�򟆶O7$<�it+�N��1~���I��2��2o�X����[�%� `�a����(�-1D�W�;�Kɴ/����ƯY���������J�@��2��$�ï�G*�(q��=��ٯ��g��?�׳iK�:'��`L�3d�Gn��v�6e����rmh�� -��i|9嶼͜�Ω�qu�F̺$ꮖ�"o����������hZw��tlV�D���{Ͽ�?��ͻNZR���_��!cq�5B�G�-2'�y: /��r묹���w�>C�W����LW����ˢ_	�e3\*n�����g?
im�/2A©g^����8N��iK�ծ�_��ćU�H 6d��#ݞ�T3NZ�b�C�_c$�X����toMRC�Q��{�����&h�Y~F9m�jw�]���Ͳ_�'_%bR��l:�Ӥ�M�8�.��N��ꮯ>i3up�C�����lӳ��J�}J%�9$c������?�@�Xk�㶓B3\�S<�OU���t
��������4�4l��w��I��X��Ĝ��6�-C<p<�8C��0��C�����P���y������&��#�j���jԼ�����:�QĆ�x�jn����^�]�� }�f���y�(v�N�D�K7t�~GO�����o��ԯ'�WO��e�,+}�53����nc��w�G�.Y8��yk������3���>3���Be����ظ���8A����R�?rH�za�E1����#g!�H#��q��|�D̫۠2�͵�C��oj��S�Y�,Թ��@8�nŜOS9�M!QWJ��(O��i(��7��;�_t�*1��S	�o���\j_���R�3Q`g��VT}�ў=��fޅ��Yp��:ب�7K&�B��!�h��ʯ�)[Q��C�i<��W��_)	1��ߝ�K��|܆��m���H���,��Gk�J�瞢��<Q�{	�L{M�>}VB}C38	��F��]q6'�El�En�3��?�S�a��=!�?%��_��4В�l��ض���Q y͡jK�h��n  Zcq6li۾Pk�K���^>��ᙧ��1kq�;�Z���8��aSwIc��OZ��N�ކg�W4���|������Ž�?@e�VL��'#�1����/��dU���g�)q�-jCOl�Q�nh;Uo�q�F��T"����s��n
����ٴ�晬Fj�$ݎ.P����"g7����6�+^̨2{<����s��I :��f�$A�d�*\>�/�[�T�d���4�^�'��v�����r�_�d�V�R�T!�]��{wO����4����?���-�L*$i�f��4�N�>A�j�*U#�Ȍ�D�@
2]�tv��e�\�ũ��亘P�EJQn��/ճ�K����)2���J�pA�έb��vZ�ɱO�`���fJa�=H��4�/��ָ�7V^4��P�]G�&�M�
U%����#��G����=N\#����N��*`�Č��_$��1Z�@V�R��;!���@lAQ�R�ٵ�tW����z�M�P����C��W�}�eK	�8ɫxW�@`E���2p�4��m�6T�j�f�%���X���䬲2��FɁK�/�G��̖L������?8���[ӰY���hwƺT��Rń��R�[˼z��C��?^�^�R�P��j�O�	����x���*y�,Sz�l�KW����j��"��yE��������rP�kD����Y���z���k��:/!�"�U�Ze�[�w=������:M��Lfm2���`:�3� i�q4ӎ�¹���a�>B��B��g< �(�y5��E��$M�o����/A_�����Ļ�$6��J�����z%^��v����e���\&��Jތ܃3������l�Yy?:}յ��08�w�U�݋�ɫ��f�o�o���w�5]��,�_M�D���5�:7�r�"������4��}��.);&�V���x��"����㴑�| !C�_�>�ո�����?�/��`��~��j�"���y+����9�U>�D���Oe��O�_�/�;kP�2�f��Y1j�R�4��{��*A�"6���A��NST�U�_z��o�60�^��L[7c��ϲ}D���k��s#��R�$���Yg�ꋮL��\�?�xx��᫱�V�}��I鈈������F6�7y�^�J��kM�,�t���O�l�M��~v˒�Y���m�^�a2�砰Vݩ�����V�h�X���o�+�8��@�|c�Cc�O��ý�u
�ǗI�˟V�������XlPJU%6&�NC�SԜ#L`�CM'�䫫�e�^v�o�lE�K�U����7�����������'7���\o�L\��0�xT�X��	Emk=�>o��aF� K�Wf%��0?���@I�Q�Ԏ��ui��K�'[zRV�><Y$�Y-	��y��F�~�+#���C)���z.�UO��ۢG�u�D-��C��y�N9G����'������N�&��"Y˸�
��X3N��������TP�:�E�]�4fa��w.z�'�}7�;|���(���z0j�t�'�����Q�57ۿ�1Q�(��=��ף�Ұ_j��ʿ'#A�#�E�M��(�=�	��X-d[yB��u�̀�.c�Yn�����}����G�'��*�����C)�Ib�	�~�w��,�C'��;99W�%7����� 5� ���vO�o.%�!k�gT��m�iV����-U#�g���fԟ�ݟHZ����=2#[�l��Ì�k���d�����Rw]��R�"z�{�	�ǣ���h����b�kKζt��(����2���p�F^�H�v��=iA[5c�y1�Z\W���J}�ii4$(bSBGU��!MN�`�;�ݘ�(�8�ߤ��Y�G<��T�V��^�(��v��7k�\�s(m�H��횉���}.3�DV��M&'\G��DAA�J�a����#�ߝj��������(����6+�M���Dݧ9`6�Z�G��k'@!������]��Lѕ�������Sb[j��P1zJ��p�Ry�,>;�^����u* ���ҭșJ��Vv��(B�̚�J�����^����mHq�S���I�S�\1�.<������oW�D��T�/`bN^Y_�_�����AFB�뤐�:�N�Ý��l�X*�et�&s���_����NDPDtX�Ҫrze}���V%|d�F�����F�� ���]Ґ��lLvA1��]���h�F8@�
��%g��PX�,Rps���kw��\�M*�f�na|A�9�6Q1��`��������W��H<�/G�ႃvIb��;?�}�!e�vI�B��Hu��[��Y.���r�?L[�)K �W&H�J��5������h)c���n����>�����+���=V�UQ�7x&�n���P;p����ͩD9||��%YL�a�JS�@vLq�Z��<�5nj��EXZ�?3 #�L?̛W�~S�6�Z7y/.;��n9aqe���m�� ��|nF���;q�T@.o�("� Ըy8��R�a.󖯡͍ț+u?���xG�x=�A��f��͞i��ڋ����y`���1{%��&���@־��U�;Ly��z)q(����D��Ŏ=�_=�L�<w��J�ֿ�Y�`{c�=O�T���+�4���g�;u���Z����ʢ3��o%�z���\�ҿ�*5![�t�a�Gx'j��E��C>^E�M:S��/��5+�b�c��>�th.J�?Z8����tǺrUlK��}�U��/Ϧ�҈�\r���(�Y���m�罇_��*�Бsv^B%��~���E��J!p�D��y7H䓝����Rv�B=+!5e��E�~I���=�.w��Pw��RoV���w�XσxYPw0�n��Ҁ�\�=�ǐmێ�]ꐤX@P�͟��1dx�1�;�o���>(^��ޤZM���l��K�?H��L��Ծk�^x������	�����֟�^�	џR
���ҧ]XwO(L�oK=���f@2�|n��8Tx���h���@y*3Ko�����<|5*���qK���!��xpVH������M]3�sB͖:~��4C��.�M<�0�����m�J}-���� ϲ��Ƕ��]V�-&lΚ���J}��jr�6:�Pd#<[,��Nw�$,�ٮt4�������"�'o�?���5N7���_���F�V���ddf�$���#���"XWި��KQM����>ħ�X��<g���å�zo95��䎢�k�����
'L�J�6Տ4#
�ܷ%L�	���aU����}]��"Qe�\���x�$�>����,$A�?�0,B6g���+�v���q6�rVPCK��4OK5̺ە���o�FH�n'���
Ri�.f*��E2�i�߱t�p��}w̳�ޡ��Tǿ�d\��,�s0{��*���Av�w�Sx�=��ڻ�	S�����e}��U5Az��%Cg9�|T+��'�6�!�6�"��n���8�h��sR�G�ɫ=�αa)eԛ/�4�|��!?�m���S��~�J�Z_
���T;�
���Z\�Ѣ]�&ס3	�k�4KS:6��ZZ��n��� w���*�M��E��i�W�_�i��p�+f�eG�x�:�7~��Ս�L��F�_���;�`zE� v-�H�O����Z%6A
�e�N>��x�XPdU�D�W$۞�t$��ţ]B��ol�D��M�!}�R�WD����!�1�>�	@���W�����	��pY�u+�>!@��;�YH���d�s��"�C���c:�	 �Z(��I`~�o�L��p�Y�t���y���<auƚ�LkQ'�$���K�H���q�̝��NNEq��i�7�s�7�y�
罴/[�.<5�~����p{(�ْ3�AEQXm+��h�0t��p�%��&���g�Ɯ�n��z:����A�n��,���ND���s�U1��2%�ë�"��ʱ�縴��xw|���@�#e6�c��Ξ=ݻ�3�ځ�/\[?֧��|�kL�ZZ�t�8�>Z�
mu�?�ǌ����s
�1�ɰk�<$�$��L*o�@㻫J~B8�ε	?�/G��ȟ|`���3�7�9Y͹�{�{H~7�)S��E��H���4��HB�-����o�_4���U%*d��}B#´\��i�FQG�j;�뀹$�͛�f���ze���[���0o��Fw^�ٝ��M���)���ۉm&��2bee��%�Wu�}��O�B+1��>{�z�7#�XŻb�4���&w�B��Dy͜��(�6���ew�u^��<e)%�u"���iK�k嗩�[k�3�k�u��*�������"�W.�=��t�lL��Ƌ�(��%�BQ�'��1��l�2J���x����7�Γ�֝�fv��%��OGm�>��}��m��	OYk�}=��]	�gs�:B:���q^����x��T���:�M���Ç�[��&�����x1��y��7��K' 5�@�!�u'5��u� `S�����r�!Q4�ٮ�z���g��D�G޷],ѷ�����+�h�+W�:��ɩo������Ͻ%99XU�YҖ�x���5`�i���ϩ"���*b���Q�vǤs��t�L��@���'�w.l/�a��C�����MbX���x��g���� }kK�-H����0C��D{Վ9��������5�JtfCp~���vo��'j/K���t00�H�F�=DuR�U��\�*R��R���?��E��N��5o�[e���a�Q-�4�EW�(b�b�fՙF���8b��%��9�k8 �$�������N1���k(4bq#˪��=Z�W�m�1a�)������l�+��tUM�l.7���k/_�#⟽F���'�[�K�6�2"M��P�;۳n���8�~�bM �j�8���)���T�
��w���a��A.���b���������?�vw�{I��g�|��k%-8/#�ni���s�uH�ҁ��XX���Ե_���>2w�A��n2�>p�D��ǜy"A~�vX���w��Ч�d=���m{��w��C;A䵕�߂ǯ�����wx��GA�Q���g�u����s�@F�qy��!����.	���_+�|�	ը�������:
k!���
Lf�Ḝ�޷����`�ə*�ϡu!���@�`�P��ᆻ�p��B���u��"]��\A��0���盉��o���?�|Q{d45e�ǅ�_޿U�*^ӽ�р�W]kc@��pCg:f0W����#�NH��A�\�G����>�h��y��L�� ��<m̌���4�eM��sC�m�%���y,�M�OU	x�M���]��G�ez�`��8W��%��3�G��e�^�+sN&qR�7[�P0?,�.T|�����m��G�mr��v���q�m3�j�~�-��ѿ��P�y#�W�=*��[6�g�}��i`��L�E�kYV����X������<�[bd�.�-�ۼ3ѷӒ���8�������ԊlZp
�$1c�_���4!���Й�6�S߼�j�sR���A�BnA���l�W�dS����`Q$7�"���l�e�qy"�,��C�-���zs��x~���B}z�I��"j�'k[}�.Pp{Mx��I�s�ʫw�'߬v'�\����a"�2,�-:<���=-'��T@=h��%��8�s��l����ŋ�=A�Uv�}u����ەx��:���3����	/�D?[3��&1��Zt��Q�;4��F�i�E���.
v�' ��pR�k�9)/���5�c�,�t�i��∟E
�5�*xZ�f��Ԩ$��E=���$�Gع{ǿ�
�cB�U��u�� ���� ��B�ZC"��%����m���K���<�� ғ���ٝ
6f���W ���ܢ�W��^���>�َe�>�PK_Q��Z^
 4���ʭ7��p����'�j�m�CVb�N(ʼ�Թ��<�c���3,��g�Q{%�T�Ϫ�z٨���Q���h�{�=���[�И�b}�����U�#7^���ѐ��R�����ZCWsXA"ٓ���6������Q2�rO9v��e��l$����Ǚ�ɰYe���{luο��2WP�o]��F��<,�+�mĕ�s^_�Đ_b-(�m�a�����`9��z�-kM���Q��C;�{
{�	v+��VF��VS*'����(L)�60~���q�Ex�B���L+��OXΈ�y�?�+�F��_��
�������,`��y �a���(���Ulj�I��a*u4��eV���-�$t�y��ej|�f��L�n�2�eG?��K�pt+/�'�f&���/i�`
�Ȧ�V�0xr�휭��J��Ð���wFQ/�[��#ɣ�9߈���,�)(��yqE���I���t	���9�[�IVJ�Y[U������*�x���7�fϕ����描���_o��o{)5��h8wԓ�I���*��WF���)ߊ\��٪}�
6t���?�?�?��g�_V�lz��ݲ��--./:�ܯ�\����"�A�c��`-��ֻ��#��k��N�V=0>�6��2d�<w�CH-���b�"-EU�N�*�*n����U�67lSSV����/*~EKYL���e��u�͡�,�Q�|���~����/1�C};��,����M��v�����$���=�������aV����T��BV��S+G�HG�b�z��� TJ���?���[�X�3����76��l������~����o�]�'HC[�G�C���7l���^b�g\Ժ�c���k\7��� �&�á���01�~x��#uхȈ��H��!���t�q�h=����DJ�0����!�� t�p]�E lͿ���l����=�պ��"���@���i��/�H�[ޛ�xa�B�?�F�&U���s�9�a����ƲW9�`݇*9�*�IBʹ�W��O˙ͻ������ވ��t��5��Rq/m^";-]m�|���Xe1>Z}Tp2	�h�;�O+g9r̼1��Z���j�ZfK�� ��t�X��`&ܘ����a�d��?�)&L93)�h���̬�&�X5����#�Dq{'7�Wg��S��6H�ǰ*
;��/��!����[E'ܵ�*�|{0����p�ӥ��a�>�x�{��9�P�0��,L�uA"�|���T��t�=�V_5���� o�({!E9��~sj>jYԚ6�h�J�W�g���D9�"ߵ�������ڙ,�*ǶM��	�g8bܱujL�*9�P�� .�9�fs���R��.d���N�fi��`nl��)}ǟ!Ƕ������i���g�l�!V�,���:#�P����Ȯ�ڱ���Ɣ;!_�կ�p�ɶ��k�CONw���[�.:��œ�EV��]��ب���!����l�@, B������������	s5���"�L�w`,V�i�a�gg_ˣf�RzD���$�Qh.�]�����my��q�g؅����
��H��_Ɋ)��Zvg3��	N)��ο]�=�0a�[�~K��=&\�o{PWɺګ2�d�y��;&�������c����½}��VWxG��U$ެ�)\6'�>��j�6c.���i�n*˷�Yh��J/�٦B5��Ϟ(;|�mǁw�(Q^-t��6�]MdC8��Dx8I�w�[`���?�5G�*�k�'����iq��������$v�2u��I��[�n^��^��?Z\6��v3]:�#ފ���lU7�O��9�>�a\	��3�UK� �{RӔn���������l�N>6؎����.)�R�[��5�G��ni�`��rH��z�i�\`5��g8~�E�u����y�#2�R��5��9��6���8�z�u��u�>Rz7����.hV<����W�M�%�{���B4=Aۺ��ւm�Z(��=�^�>��"D奎׎���1Ҫ�@�P�X�y�g?F�ŨRh��k%����>Sv0#�I�37=�r�������݌��2��նȼ"�4\G]Ϲ���z:C|��W�Vc��U,O������%��N�j"�6�((���r�7X^|������
G��O,�_�<,q3�2iC�c��߀��<���ٲ��ƽ�-Y����mC���G"3r���a��2c��#Zus�h2����|�:��L(�j�'�M��)���Τ{���a�4'�� D��C��l��.Q���a i� 3Gr_�Q����Zd���^b������9�q%ah'��ʙ�B�^.���N��Hf*ԍť���:Cz���G���>ɯB�[cQ��Py���?���P)ѓ���'u��oK:���0~���)E��
�:'�=[��hd��@u4���}������5���g�}����^�a��TA-HX�%t�ƻh���56?�-2J�J����x4���T��_�F
��4��� c�q�_��.��*d�.��b�/L��2t��u˛̱h���D�p�qd�D&ϛ��f�&}b�o�Ą��| $����
�U�K�|��d�v��ٹd������;���׆�'o�:�Q�#��4Rc2H� ��z�%�Iŷ�YY�R����G��Ã�#x�Pk���C�����0{�/>���9�������5]�$�$_W��{;~�Ggqﾸ���hI�j�hD�̿�A���E�I����(�7�L�:}|�L�e�8Ѭ�3g�UY+������-����b�uz�_sb��;����γ� �X� ;Ҳ�/�M�W�_�*\2���ކ���~:n�����]Q�HY6?���O��>�����߉�v��-�7Q�x��¨�Z��Fՠ=�@=0�V
Z'Q%s7Օ��M��y�s�iI��x֭�Ev
+�3%8��ojKٹ6�xc,��K��cä����0����_rE_J처���h����L�Ir�i��z�V��j4k}�D��I��;��wbq��>�"�Ά��٨��4l�lb��M��9\Z�ɠ�l���Fh-�o��N6� �%��O�`Do���~�<�J-\?����(����ʉ��n��$��8�\��uK$�<��!c/�X<7)�/�<"^�y5k��g9�kgph�
����Gu*�8��j�ڶ�͹Y��T�H�5^j�K���*b�w�uf{o>�;��oN�jG�G��T�C\\f0�nxn�}�Ɏw)��o	Ox��M�I��u�r��>��k��6�N݊����&8?
�*8���<�C2J`�
{铰$,����]���H�ӡ�� �2-��o�!�?���H��;�I����ͨ�̴�'�;^��k���V��+��mZ�t3���/����t�� �E�R�K3f�j���_�I����c�7��եo"&�W���dx�A����۝��?���Qjrv�|��V[y�neW$6/�ˡ$5�?q٧rK?l$�����;��g�Vu�x����nd*�Mo��&��50�V`���l�jd�pHֱ��b�l�o��]&�����Lz��EEgPf�e�#/�t4DTAB��x
B��-�o@�7`ֳ'�B�Y!��7A��R��,9r�q�H��!���\�@�|D~���9v�Y]��t�]}.d�®z)/J�7��[�?%�>R�-�x�F87�}�X�k���~�0�����\���b���:A���|��2`X�hRh�N_q�BH"R�؇�0�,<r�wIr�kB���_��0��Z�]��d�6���=���	��|��2��p��rQ�-$��HS�	��� ��o��c�1`А9Q�4YH+�)Jr�ge$t�"��q���Z�y-�HUe�'�%��O�	�À6�1�tG���'u�V����>��\����ڰ���	�+���K��B��������EY����X����ZAQ����cТ%�Y���w֡ ���W�C��7�8%y��%�V�����MU�{��N�	��������$2�7����ޯ�,~�dC�歭��\�St(�Ҽ@umn��7�'t��_���|ˋ<B]���t������D�����&YF;��%����v��t����ш!I;��WNZ�������2E��9"mTkqf��R��2�'�'�����Z߹�����tp�\>��2�=��:��Z=�/��F���u��Q�k�GOQ��0�7�X֮)���F��܆�J��B��Ν-̎�sLY��Ug�W�$����X����c��Q���>�A��a6�����
�@m\�&�P/v*f`$y��"�
����5�_�lay=x�4�����1_o�����mư��9�1 �+m� ���[{Or��t����W2vX�g�jy��%�y�:�:���'-��p?14N[���*�F_�2����o���FZBJvӶ����<�	m����,��E�k=RBi��>Ү�6u�t���Y�1��a�ş~��M3��ID}�Ŝ���I>��U���%A��?�"���+5k�W81q[�����"_����nׁR{�H㻹`:	�@�Ѭ���o���W�j|�"eI>d'c��o}b���J��֨?���y�-���@g��t�3b�	z���ԡ-�/)I��QP������]�����`6�!9�����y�W7MG��r���"lZ��R�R��l�iVwbV�;炥���P�o��U;�&{>��cTtx�8JW��F�Cp_��& ���]����Ux�������Λ�	���b
қ��@����.>�m��y��8HJ_1%��/�k6l�2m�Ѧ�R︵��a�9�|�e�2f�G6�"b��������_�9�=��[�$K�zj��^9�M�T	l߿���K��9�b"��}[����|Y���#�pA"�A��9����|��@�T}�K��#"���Z);J�?JVT7�ػڢv��Ѐ��m��q��-Π'P��}�@K�Fŷ�rt�o�ļ�	��e{6�뷮�z�zշ[�ϳ�s�8��c�w6���q�Q���$��<�G�u��c�ѫ��!�>�.����O�|Ҙ��ә��{V���S,s��::˵�g7q�)`J_��Ħ�uO}�3��iyڜŇ)zde�%5�Y�A��u��M�j]$\ñ�4�����p}�Z/���7�w�x��)r�[����t>R������w2)_����W��� n:h4~��rV��=Aq����P�sz΁�~3����o�vCXu����v؄0�fjoKl׿w[�xm�"��EVJ�o�a`�	t!΅P��D�_Ώ{�*�B�=<s8�W�����7S���]�!S.�����S��f�BO�N���I�,Yaj��0wy���)g-@H���Wb��k��p�ˠ��#|*���ׯ-A�Tq�&�>�9����11C�i�ͨ�����Ϸ�)#Z��)D���v�y ���Z���~�J��K8��R�6��� ��f���s�FW@OB��9�T|P� P�1�Y��&]���e��̡�-?��5��Y�������E�}���<̍6$-��E��C�����<m���_@��t*���vB��qH�%:$���X���%���i�Ʈ��?!��c�~r��c�W!\H�2��#�mu4d^��L�=��wjXRùrJ�b��7I80�����"�]��S0�w��@����پ��>������3�Oг��8w�'b��;�j3�:��Z�9�A��4�Nх<zˈ�x<��)���Ue���p�!�����]I�� �p���x�(��Xo^����	ɴ�?T}w\�KЮ���#�DQDAAz�QzB�R�7�$�(�4B�&��^B	$�ޤ�J萄	I���w���ewg��y���}��䢛��[t�.N�I�Wx�gP�f��n@@�"�z�Ů.�wo�0����$�u+]��򛚣�Y��8Gbz������2������u�����kG��%}��m9w蚓��OЮ�E�w�������EG�-6�a�N�%�1�\)��q&˲ɕ�K��@�����Q�h����+���XǭL�H����`��뭔������cHO����e�%5�,��-}��1�i¢s�͉�;^o��L�Ӣ��׀e���\�#H�7'�z����ނ?�,����FMak�ҺD��~4iG9"M�A0aP�A�4{��]��i�X���Tg���.?����s���
*�X\��%ԎR�$s���U-��B���Ǳ���/���"7'�z�0��+��RL>�׹�s��.�)p��x��9-�h7FȑBZ��k�[�d5�MRG\������ˁ%. /m�0�Ï-�,ΠEN�wZ�oH5<����6͓T:?�:lé�Rc ��4�����7�}=�g��SV+��K^�L�n/��ϵ��{����=+G�������WR,ys��c�TuO�E,�r-e�����������q(";R��w{*�C��׽g���+	UQ&=�eĈ��fŦ��ύ�����_�������V�l���Q�-�p�̀d�pr�4�q͚�k<�N͗�2=h�t�g�~U����-eo���y_����fJ�q��	ǗU�������EM��ɼG5��I��dc����=�R3��Z�Jc��J�����u��%M@O�8��f�U@#γ�>�c6�ok��v�k�������x#�u�Aڨ�>�W\���FR\c:p��ä�W��"�s�ӝ�Q�Qd����HL f��@aw��"�1@��Ua���ʦ��&5�|�)~����"\�7�YC!�w}x������������w��9�v����I�[5C�җ8�|�T��K\tb ��}��cqhK��-\�dbF�Z�2$�&&}�u� 6Qw����'Ԅ�_h�
X#�>�٢��]�O�"ҸLM���O�����<���g��b����_�r��TI�.Ǡw��V�/U��<\�[#��T�Z��(��e����K�������ĵ8'©�g�ա�U*\�\m$�2%��`��0\��9�}��S�!���3F>�ss���sZ�@��Y�|�X@���A�����,@��e��g�������_mt��\5���2��'�ȏRof��fq4����4�������)֯�C������殹�{<�{�<6��N����y���ہML���>˷�cQ��0W���AY��|��O���m���>�!����d�#���x��E��d��|���ާ0e@�V[:�J�Y�P\��)�tg��?�՜�r�$��}p����.�)����L�J��K�!3e�lV�.�17D���:'�LJ������A[�t�r��s�b__��G$YǷ6�R�x�pݩ�<�7��V�Ռ�$%�R.q��*��X�_鴥m�;���#�ss�X�X�W���1u�o����A��r~{f!�Y�0]�����>7�,�#��c��(�o6�J�C�Zh�]��Ɍ~ڽ�~{ y�tR2{a�U��]{$�����[�I����Ľ�2.���:|���<�)7cb덀��ID��o���7߄W=*�B��6����6�jk����@�P�s?b��/��"�]e8���V�@��.�fb���W~%��3K�=��ɥ�I<���'w���l����O9īӆ�D�/��8�A+?��ҽ��h������3�'��-�|Q���q$��CEI�݅���l��&���f�@�O�9�}��_1�\c>_w=p��2�����4a����Uh���ެ�ƁNG Y�k]�^��rm��SA�_5�Q�actfdK53����A@t�6��</PC)�v4�,\`,=P�����hF�(R�3R���,�.|��X�<׽K:(4���)�K,H	��h�w�FB�V=����(��wVW�E��Ǣ ���U�X��L�����U5n�A�}D���俫h �����%���f��4�ݞ�o�M�l�*i�4c���5f ���aYK�iD���`���g�����*3y����KJ ���E�j��crײ��8��� tWA��*��;T�R9�yO�o��[�g��;�n������7T�b(o�{�p�,��n{׍����o	�R2���M�=���2���e M����2��y��Ƞ�7h7ˊMr�JҢwWO��j�vd���>� ]�L�i�N�|�]XYZ����8�J�)	7}�$a۞������\��p5����A��`��ӂ�\��^[ANv��	��0 � ��HM����?�`xz˞�_DB�H��u�
�{�'��+z+�c׵�H�O�4�2�;R{8.�5���~���}oy��kt}���$���uh�:i+��V�(�vxUQ��
���]Pbؿ
����H.M�5���D��4u���̴?u"-�M�C�1��7��OB�\B�a�21,�T��sb���U�y��d�7aҿB���ּ'.;�a����|��%&���\8YqD�/e���Kjl}�@~��^��>�h�p��D]n�;����#NdC�'9ޘ�l�w��J�.K/Z�1W����?����7�%R��Vۙ}]�����fs�sx�lLۣX�X�/-ߩ���֍J�-H��_��` <>D!2�3�v7�M����'�$v^Dn�g��iuA�h�e��8��Q��.8�u��`�~fo�ܿޅ�N�v��VN�;-�&�>pG��|�n�S�ʣ��8��#�遗��������f�֣s��яR��y�X�#-� �"a��@?��I>�?�_�XG��L�5��++/����y�n�����������ݷ��l��`�7����t?�l����J<���*���S:�.˫�=8���TԠ�}g�5��}�E���	^/BUT�N{�3rF�q�j��g����/��K]����Q]K��������歩Ƌ?y�b����ɥi��{VG�#�������P���;x�\��#`q���Ѻ�XLĹ����Ļ)�ӟ�;������}.�����~ ��G�-���$���芳�~�~�PD����2�ݩ/y	��9�Mh\_n���B:�T�f�8�P�]]�Ѭ��j����耕�i�.��7Ic��V����L�4�+}����Z����fR�L�z�Tۚ�q-�S��2w�"=j�`�y���zm`�aZ�ИF{(��`T��W�%�RK.I���9��]��Vóu{2��m>�n��\-ĥ13�R*ҿ�[�
��xY��O���ޭ�Em��If���	���*�i���y�� r��^�[`8�ʣf"�Z�~�}�[�"������w�����{��\x��ܖی����oFSK�����%q dQDAIH4����6�Ney��ӣnQ,"�l�罻z�Zfv�nMh1Y�Y�����E��/5p��>�+-<M BHk�_:�Qf�:��N����c�����7�7e�Fq���-Nƒ���w\��� �.�.�{D�, ���$�����˒�S=U~�#k�T\p+�M�["]��
�����+{��/��e)��R��\8]��J��C�QL�=l���U���#`x5�4�-���ҭ�fs~K�k��7h{�,f��bǡ��W�><ё���n��9,*W�)�7�`�W��X72�p��4�=�.-@`�I�&�J4�l��	9��k(\\5Il�^3�B�[)Z=襗.�����i	+��-�uJ����w%~(08�yq)���Ki����ѿ� �ɉ�����"g6�m,ID2>���7�|�6RYk"8%�Ĩ��X�y��n�oR��}�!����im����ǌ,��:�t��ٜ��3�W�ݒ;����S��s�4J�ٛ�L- ���]�v>��P��H��t*�.z+h�M�NG�Ub; �(Ƌ�xR��vl��rdZ�7RH��/ۏ%N~��($6wjT��@o���	��>�!�1���h!�Y��������A�:o��g���["�/�Kg�nM%v���fڵ�������׭	^�,+-:~�����{�ۃ�݌��	�i߇n0�7�8IN�G��OHG�z�4�aW�����1��i�;�y� �e�s��ۍ5��䠧z������`d���Ë`۵��_���s\얒J�V��2��U�J=0��OT;���ħa�~�Hx�_����7NA-������xN5zQ��+B�Y��OT��t�✵`̈���ߐuuVU��j�1�g�(>n�~�MP�n���]�K�L��aVz��]��%�/�q�޻'�G��5�� �e�6��rc�7��0X�Fmhl�%���I���������b���~������ɑ�9�U��^�v��q�N�O��*���(�]c�l����w��̬��6�,��T��lN��J�LM.���M3�ʕz��a\\]��Ъ?,#��[s<~D/����O��$�P`��6���I��`�?o�N�\��^���5�%m��[���bC�� 	��˫��w�:d�?��k�v�lv������@���J�R�lG_dQɑ����i�,F��%�2Bʏ�K���z������fd?@�'F�v��wB��-Y��q�SeK-E�r.KET��}H+3���'~_�X����!�~�i���yq��.�����I�F�G�V��狟{:ГU\��&�ν
#դ8�*�{��t���L&=�&	y��z<���e#�;���諾�o��8)���Xu�����$�m"t���A�Z�&�-/r5񥩽��S���"�5��tACG��Y������R�.��Bz��/�":μDPp�qH��c��1H��tؕ',��(M��l���}��rv������
�Ss�����^�O�u~�i��	u	���eD�i����r��wL䱰K��+^>s���������m����*�)�|��9��n&{zv���(���;���2���OF�@/��i|>��NP��-��4���C�ov�+&|
������u��ɲa��v���je0�F0������c6�{����5rr�Zv�z���[�.A+�ή��U�o�k������|�i$ {��!��Wջ"�	��b��M1��xl������떙!
�wõ�Kq(�؊>�S���e�A��K{sb]�d�����Wu�j�����B��#5 ���hr���9���v������x:%���{�>��i��Ƅ΄���h!�u��+�5�n�ć�b�;3"(�"z�k�[��6.l�Y�N�ąF67j���֤b�t:�6m;
qܦ����wY�v<.�#j*=�v>a*娣������+z����|��I�����uӏ�sEpћ�xl��وhȫ��CpP���K��fe�ɔ�k{�
�`b~��ܔ���V$��LfU.��*���bs���47�~cH�?�M�$(�-9��"t��W�Q!�ﴍ�-�����#�%,��\��������QTԴ0
	�f8Ua����8�:��R1[���o�&�gk� ��0bN��d�)�:�YvCsCJ�X�ٶ܆��	��.�����7t��A@,��k��d�.�I�&�t����e��/���$K�a0x���J�� �X8�Z�L�}��X�i$&MVb���Yg]�@��|V�TR^�k�[��j�Y��p��z�g�H�*	���_�h���RF�MvVm���%�~R0e7�0B�S�>^��3撧�Fx��i̛v���frw��Cl�&�y�{��N-�'��Ey<�X�G���%��㰺{R���f�`$�v���F�2#6e�|�6< C}�(ױDx����\�)�#�9Z*�E:d��>�o�:�B���P%2�3�%~�}u�o�K�N����3���iV`��U���	7�-��L�t5����04��w١pU����M8�-v�7���?��H��ڷ������D2�3�ҭ	��Z6>�ݼ�"\�N����=�/\�"���Y��@~��������lgsw��&h�7~�(�;���kp�{h�O��Ӎ�RDT����&�i���k1`ʷ����A��(�NNs��/�ٰ��N���e��#0ZS#[׀�6����Zh��my���7\�(��(�M�i�QP[Oq�2��GPs0�-rY(�C�o �5jd43Q��oǌ��";�%G��"��<�L���o��q�pŋ�w������̈'�����u#��iY��G�}�S��91㋱c)G�{qP~�%��T)E�e0�%���y�4pʢk�d��F�.��ڽ����&Y&%��B�2/,���N&çj��a2��h�c�P�ڙ\�a�E�}�X�<^��ۛ�L�a�b_ �8��b�;{�G/��/�i
��%���oE�.k�R�uiTNo9D�\�s2i|�B\kD��v�Df"K�~u��CĊ���Ы��*b=��v�iB�:���iv��kT�쬑��[�6"����Й����%�zٰřn�@��?M<�_��#9%~�*N��}���Bxzit�I��z+kM��h�7l��8���r�\�ȳo>$�J��L|�k9�(�A|[��>�f����VT�#�[��i#�/d�!F�2�b�|s:���מ�[5�Q���x���pt�1�ko�5�����K�O;睜8�5�
^�������U6>{����Q���0���,-��	R�5.�Kw���5��\�뫧'�u8��qq���vJ(_��xK��=�����G�q�t�����<6m"�%� ߟ��ǺT�2��9����w�;q�?�b�2`�!��{��8j���Gp��XsD�7�Guu�}�}7��A�y޲���ZA
2P�6p��1�X�)Z�-�~�޺���0�#H00���YI�V<�*�L75�\�����*W��"L��������v#��c�����@)x����䒟;(d�ڄ���K���S�[�mX7S�W�W��Z�s\Z}G�w������R�\ ԭ'>&ܘ�G�ď��'t䑳+7�Ւ��I�A�2 =g�z�꩚D���{۾~M�h�G�{���+�����Z\61��V�}?!G#��b��oh�gx�����a����UL�yE�R�{��9�\L���%`XW'����lR׎@��E���EQ����sPǌ�MQ�XGb��������L������'��+�4�6��r����uV:V�{;�s�6�в�	���fJe��1�޾�9?l�o�w�\d����e� �ʌI��u5io��8~���~^o���m�� �80�[�S�66�d�{�Q�bV�ublO�z��S`3�6�2gxS�6��0xP�u��V~����(/8'M	2�N2���?��^��g��]t�
� -��9�L�N�6�9��Pw�Y�+�!��~*�3Z�p:���Y��^��Y:��;:�ƴZo^�[)�`0�.�Y�����:(�>���I�������<g����]r�7ݴfF �FZlb
�μm�J��h�5�wt{�V�BQ��ݍ4�v����e����h��>{�q��>���DTPC^��U����n-�ɻ����4\�<gN��u�	ܩ�f�:q� ��c)��7��1/�r�����e�v�h�"W�+}�~�fh��1�Q��b�gt�r�m40'���9���Pw���O"�O��Z���"$���o�$tq掆�j<a���6����ۖ��_�eX�U�J�����p�����3泇Wl�����eڦ1����Y٨����x�M��\�a:��ƨ�:ܐ��;Ca:'�.���l)J�j?rI1.q�F��6�"=z��@�ٯ��	�hٖ16EZ�St��M�_ e�6�'b�4p�-%�,aR/�{�J>R�߲�5"�7\���I��̬w'>��nEJ�c#��8x�(S֊8�c�0B5=\NLl'9N�ת���
	� �\��z��g�ʚ6��.�I�����E �ӟ}����f�w����93������i�W)Z�m���x/�~����Kfʡ�kH�e�|�sjhh������;���h���լŮ	٣�.除�Ĳ����Jg�SRgz+SsR"����\�D��KK���|̄�C��2�ɚ6��3~�տ�t�L7M��_hh�4��֮�Ha&��x]�CQ�#�ޏ,k6S@�����Q�0�S8#�c�*��������vz�g�Gu�D���A�l�|}D���%'ˣ�#6U�����R�	���Q�.��&wܰ��2q|��kb��k�I#��-�;%�](~B.�c���.�����*�<e�����@��d�lxS8R�<9s7�nvp��]�H|B�r�vz�j�� ߟ�����kc_8*�s�$��3�1�E�.�=�ߖ&̵;#���p���0C��gD�����~��dޮH%�#V��)���y+4q�&�r��B�N�y��j���v�*�>�{�s�l��uԮ1���ߟu���I�
�� 9�ۋߚ4�ۣ�:�7�o�?���� ��� ���*�.�%Zɛ����2��V~7]3����>5����a�^�Y_��j���������������{�QOm���3Q���̫���''`^--�1C����C��|;�1A5mgO�(M�7�E-��JF|Я�̳Z���l6�d�	&m�[��we잓A�*�뫋�~'cI���f��Q�p�CɄ+ �Y�S��~��>��ׅ5ؽ��K�X�u��ΧR���"���#C���]�m�����)�%$����
�P)�?YY��	����b�"�m�_�G�GǏ{�s_g��j�{�G����s�2Y��78A0L�Q�5���� ���K-0�M�~*(���&��m)>��߲ �" ��R�%���-�k�`�p{�?/X��)$������T���5�c~�@�8��#R������V���Z���*n�����kÞ��������o+ܞ��	�?���f��hO ���������J��[��ϑ���R��M^
��
�Cu�Cd^���/&Īf1�K�[�y�� 6L_�Q�����R��
��1����VwS+��<1LFV�{8�}<F�����+���j����k�ܪ��M_D3�a���r���
NL-��U�,�؟ܗMa{���fS�5W�uƝ�U���(�<�h�LCd��xˎ�_5��`���D����̍��>p�h�� ��RI@�I�InD|�,?M���)F�wz��GT5�>�{��{��6�[pd�G_�R�G��̊��֟��/2)��6���D���K�M��w�����O�C��T�j��yc��s�diX� ����SYT_�&���X8v#>�6r�*�#oee���q%��f|i:j��$�⭪K_F�$� ���h��n��S����҅�^��ݍ=ٱ́E�A��q����z��Fy��d�UE!n0)*�L�I��D�*	��ŮaU�z�*#��}�zu	5��NG�yJ�(J�D4��S��E�?|��f[�{r�E6�����y�?<�!#P׼�
��=��>��`d/�	~w����VZy� $�2���c �Kӿ\���HH��ϨT���\���B�ڲ��<SƷ�%Ζ
	&/�_م�����KΈ�=���D�ǖ�xo;{ڈ����M��T	�"�7'�?�wz<��"Ɍ��X'6����G�|d��;}�q-Ɯ�a�w��k5y�6ܲ��A���Ûi�	1�)��5��)�IÔ�J��I�N�s=#x*�،���ɝ>�׌}j։��һ듦U�{[#Ԯ�D�)�I;O��R0�o��P(�8��+QH�ڦ*+1���a�޲���6WD�nWO���C�>Qf
�ߓ�3��������/
4'򹀌�Ҫ�h��?$�!�N�꺏.��KxC�n��W�M�R6��D�y>�|��Fj�R+��Sz�4��AH~���B����-t�<�=ۑ�1{��/�C̔t�(�F�ɿ��|{9Nz$����1OtoG�2n8�/���ڞ_�r �y1�|�:�UK�ZXW���Zo�N0c��l�əVg����|�����L8����L�#�k����S����W�G=��r�eJK_&�H�W��B3�F�;1>��o6��śڤ����Ό����'�����������7]�9.=&�r�K0���Q�B'��k��f/��Ӟ�)[*��p�8;S�Գ#�o�p/�x)����C�# :��5��}��|g���)�3m�A��5akp`"`*���i�T���a� �Oh�����n�$�+Ԅ�B�ix;��8���O����'��{،X��D�o���s�n'F�B���Kv�k뢟/��V�E78}�&s􋋓ʓ>H-*P�p�.�锄H��6���E�&�ۦ���AN1���>���Sc���dK�e���x������]�NG� ��^{l�N�!�v5%>�#�>ɍ���S"G0ۈ�^.υ�U�,ߐ��Ti��30Q�E� ��ef.&R�, ��u�ug@]gFN����5������*"�:�^z|5�D�DԿ��S
��|�R�F��{�dV��d����S�ƪ���5a.S�R��=�����d.�5|x�jݳ�=.qݗT����H���a��\#B�E��Z'��q�nM�
�2{�����ƪH������0�=�F���d� ��DD��؝>!;0�1eդ�+b������E^���ˠ���q篴vڤ�$�>������ǟ*ī����`aM�����c7�2������E̒�����x��햰E�X��z7������0;CY�_���rر}~�"]�-3�_����\�,\��~~���גv���Ǒa-#��H��B�a�~����h�m$��3�å��&̷VvhݶZ�,�FnO5�=݁�W���6фP;	�u�O�S!�#��ƎӼ�~��hHٽ8���F��I�����~d���'j�0�$�13�V0Գh�ա�@\ATDMT��ad��uflgn�#��l
ﰹ�,��w�C|��<��N�_����s�0����k.�;F��EOo�$T0��*�=K�����Rm�-�;a���x�F�9��3MΣi#8���\3I&��-�J� �դ��)\'���!7�"��j�k�����yR]d�JI���tf^p1
xw���\�LzhK�צ�=�w��éտ�٬X��	���,���c�J��*��jr����������#�^l�M����ɋ�%b8�-����Y���U�xVo�ho1�����*��HZ�s�F悼��$k�O~���|hg:
�y3�^��:���ώ���K\���g찡f����W��-VT6�\pޝ��gl���{�:F� >^K��o����wV=����E<jy+{2��EMK�ˬ��	�o$9�bF�,�F�>I�oe�,k�Jo���]-����&��+vu9�����6DP7�n]4u����&��*�o���:�5���_�LRpNY7~�ua�W�I��3�O�r���H�ٌ���Lp���?�ƺ�_�����
աBT��\��*dE�"��7@@B�ű�C���Z����7�L����P�,��L��G���M2 ���������[� �n��0����V7a�)$��Z:Uy�>���)��`L�� ����~_wx��R���D M���v�
���s��3O�ht�l�����v���g�3�g�9��e!��g�{y��t�n���Y[�9ҹ���Ժ�% ��>��ybް�w^�9s�X=?����@�~Y�ߟƾh�='D���H��EK\Ƽ��|51ܾ]�L`J���c�S�`�ֈ8�m�(�ac)*V`]^����+��౽.;nV�OcX����Iqx��N	��'��v����A���Ԡ?�~��دsK�u��-hK�k��iR^��5�(k}T4C1,��>0YuV�]����v#E���{��DV�ؿ�IwVf߽�ͅ/R\���ʲ���7�p�d�K1�Y�����#"��%�L���J�柣�#.�~��2�dCl��Q��KD�/�!\�ê;>��f�H��h��P�g�!y�a���]�W�|�!m�](M	����Ϣ�g��1׉�K�&��!��<#��.��&q��݈oB��5o!�x@���v�EU+�;�<X�c�����N��{cj����A�� ��nD`��C������X����<��n鋷�56��4@�ƨR0���;k3?��B1W��M���x�;�q�ݒ�X�A����\��'�R:օ��䆽
��̏�|?��WUK2��]Hl��wN<���<"���eK��K=˝��5mf_"�\����k9�9��}Gq�>�~�:�5�%0��iBjvt�����R�eդ�9�����f|{������lt^�~�_�q��T%��۷/ˎ��۬��{虰���:�B{c��m�SI��
��t�3oA6������-�ϸ��ֻ�=E��G�W�c�︹=W=��Q�>�<��T�����}�-���,���>a���W�����B�*�!I?�s�hU���a^�����+�VyM9��yof��d���^�� �+�����:�]�͏�eGs&����E���np/���.�����:��q�Oc;->5H2e)��N�5�*¸���/S��c#� 4 c�J#lo���A��A�_������������B�ʱ4C����L۝p���:�Ru�&��P����&�@�����Mo��^o�}&�ZhE��^O�R��K�$>�zeHi��ack�07$�̐F�ᕜ**kx�.�/ 1�?� ��=����^��ɡ?�7)���mݵ�C�kџ%|㒯��}���^�`(�z���aU0�̆��:�{���<�c�`��h̡KoOF*ݒ�1�6ڲsh����GM����]UQ����M���j��C?��'A��L�.�m_�$��:��o�$�Mb����ϵ,9���c�]wYX���x���[sU�up]�5J�.��ڲ�G�ᅾ�BGׅ�:N�\��5�������$���'��//d3�td��r����"�Z��Z���[���m3�r���,Qh0��y�ЅӼ:�(ٰwwD���R(���+�_h�C�.��?t��������������-˵��X51�ޤXu{f�>w�q�iC���w��5��U#!w�QW�0M	F�!p��>z�'ة��XmdJnfV�lnB7'���,��Ϗ�f1��hT)`� }-��Y�ٝ�S�jOz�BH܆����m���o��Z?,K�[K��\�Xl��D�S^��6q�U�r�=��7�-����nR��ZS�Ꝋ��1�R����,j�i�x�S:
��%��d��.�zr�S��B��F�1�7���[Gl��8GXk�L��;���/g\y��^%�"+=��A�NF!R9:���|��=���k�X���#�gϑ��=^�	;(P��!zs�8�ߕ���NY�mY��L����z%��d?4�ƻ9���a%N	�/�`(�[����&��V�)άɩ������ŝA��`2Hi�Z�����Q��:ѩ�v�?�x���H�ϡϽ6���*���D'I����v�$]Q�����s��	�]�~mH�D;�78P�F���|�w�6+^Xo�	��5�*^T4�wz�\�p���/��",�@��c��b9,#Ez�lj{N��3�_�!��y���Z��^T魌�0� ��I�U~�ʱT�qcVk���͞� ��z���H8����_g�{#��ٴ^�oQ3e�*�maI�%0J������9�v�����)��ו���̎�Bp����c��; �`��'��M}�y����O���{�
Ń�'�����Gv<W�d��S=7��	6�H��K�/��@w_��L��c��u������[O�X�c�~aC7VC��
'��̥�^������[7�Q�(5ƻ�s��/廱R�����N�{��3���׎��$��B�N�]���F�z����KuI�Vtt)�\I&���6�0x���i,=���GV	�y��ߎFho�Y��(6�N6^�/�{��d�چ1�0����&:�߶XWc��7�{G���%��ko��p9T��O���X{���~�M<e��(u�ȕ\����%:{K��:$� Z���}��/s�{?�ɗ���(�y���� ��wk�gg��ox����N�g�Wӿh���rWjc�k)�<�id>ѩg���^����)W��m���/�B�i^Dۢ�Q�n;g�?�?v�gK�jBwj�3j9w@14p��:�pf5�Xx�]��S ���N�h�9���4\��V���@n0|4�n��up	Xi�Y�o�(Q�Kؐ�5��y�5�*S��)��	��=b�)q��B��� �����F)����M�1��-$��z5vd�\���d,�Wl~�'�7��� �:s�%B����?U�YǸ*#�I�f^�{)�/B0��K}�v9_V���sn<'8�l��%����|{3Pkސp�N������������r��::6L�O
_��?�C5<Rح�X�Ȝi�0 j�G����Ĭ���l�9�VL	�t�Ww��n�����	��5����'�F- �!u�;
��?ah͔��P����CQ,�ؙ׳�;�ѻ*�S��0>��]��ՠ{�T�+�;�}�Un,�LM��2'�K�����
(��L����]B%���Q��E��ٟ/��e+�\� �k=�iE�^��R)�qT�v�1X����8�����.����q�厯�ܝ��1���`�t���h�Adxs��rl�'���׬�Oo�#���]�fQO�u	�]�b,��꒶b�Me�~*��?O�ܜ�s �T�>��]���
��_U��3�Y���|�k���#�/z7�9� E�����R �Q_���@/�fE�"~n��0sR��^zQ��z������4�YR��Hиj����Z�W�����4��V��{)%ѝ�O0/�3y�A9�Jxy�n�״%����J���AS^v�P���w��j6�U�N6����*��/շ��c��_��'dK���퐫2�&�8�y��I�����?���-���mg�U������ң��p�ȝ�)�1N�Gּ�+�j�;��&^�wW/�G�e���o�|��4@�F��[,.��𗸤Oz�/�Os�C�Y����Z��r9j,dY�p8�'�k��;���H��H����$��^�ţ�S��l�:� {'v��<���jK�[1���2/h�}uͷ-��'�/G�oK�Ĥ�-���͒����U#�'�yyG�'�Z����^�q����M�N;G_����\��jCl�K�|�Ri�
�����y|.c�'��8�M{h _^�TZ�݆F���N��<�l��	W��r��	���vk[�u�O��&x��I&���uZ������<�r�H�D�e��qGq��c��J����w��{�b��i�&᫪�E6�Z�����u�K�fa���m��bæ�ł�1���u������Og�2"�~Sa�n�>�#�K�d�QL�@�;j`��[���T�x���<�nӯ���«��}��5�h����+�����l�Vn�0�5m�G�jw+�D��E7�/h�/Q�ʹ������#&g�(����釒�5��H��`2�C�z�_�;�AC�\��9ѬY���Ѡ�y%ɥu�3�7l��냯�������e1�X���`"D����4���1!���S�'/�'z��7Mj��5s�+�z> �y�{��ݹ�;�BB��*�Ȁ�vXΪX�#?3�A���Q�݊w�:~j:Z��;IW��ƫ��{��/�7n���ּMr�#ĂezK�bٱ��\�x��L�A�=�/��©-�H��y�_V�/��kyb�F��2��rj8�5�ve{l8���PK�)�cެ����r��(~�r����b?w+p�S�~�)����Z��O���y���v��7��Iҿu�O��aH��G-�t�#��U�鱈+{���rO�/��;6���5b]Yw����M��<�Q5����p�~��J�$wa��ãD�{��SPg��F�|k�;)����w�V���o�5���8���*ì������ve��3#xw�~I��1U������~��\���dG�}d���?*�<Y���P�W\@,�a�?_J�B*1�lem�%jt��.�3��%��G_�j�����lD��>N8���t�2�W>�_~��w����g9+jtT����{s���;,�u�&�|YJ�����C�k����F>�Tj��|��̍�s(�t����L��i��V�z��=�l��a�=�N���]�Z�"���R�I��k@�=!@�
�H  ��I��^��=�&��������*�f�3s��sϜ�$���ʑ�&N��,��|w.�Z�j����7�w�Y��l�-S��"K<�z�k��ȀPu�*�^?T��h�C�..�&�,�\��sFi�;d���k����a���N�K��"���R	�b������Dު�x]���Մ�_df��s�c�E��cI�{P��i�ּ�~�b�a��^W9X��=L���:d��0�}1�G��+��ۏ��`^�p)����0��9�G�%�'�y�V߅�\U�Ff-��(��/�h���f�5��F/k{k�%w���#�օmV����.��L� �{"|6Ϩ�s��އ�c�ˑu�p�vи�Zxrw�����sj?�6�ƴXy�(j�[�=
-P��z��"�����{N�����߮(��糇�MZR�%k���j�*|^��^�C?Owa�͂���ä����.\2�+[��+(���)V�֨a��HK�5�,��_���զ�h�����jpHl�+U�A"�=7�ۻl��y�_�N�gb?W���&BCW�^�[�0��.������`�K����n�B�q�Q���2��ޫ�_�䥱��
}���>=a�sk(���͂�Y-�i��Q���cSJ�M�Z��DXg�o0�TmN.�:��;qq�3�yi�r�>`W��|s��H���:@�����9�b�]�r��V�ua�E]�'�`��V��t51e+D�{���8�
����I��Ӳk�I��Q�A�zt�s��(愺Ԭ	�@.�nC���p����i���$K�l/��h7Ot���^`�@�^�|/�m+�٥�U�I���C�p��a"j�Յ��ϲ�H����������Qv����u�-�eC?�Rd��tl�ĥ8o7�@Mqeg (ҍ��%��4�������*3��ʮ].?�0��K+'��E�L��?�/�F
w&�Ot�]MX�(}ӻJ$��\��P�:��]d��ڊ�4��p�9T�>�@#�ܸa���!��}h=�Oջ.t)[��9���ձD������[)�P�P4���2B�g�Pg i��v�Ԯ����c���rʶ͓uֆ8q`��Q��uѥ֥^O��iٮ���;�'f�fuU##��s�.���4�S jS��Ō�3x�D��X���4D�.�W����x ��V�{C��*��m`����ԅ8�c, ��y3�u3�LS���&�*��I8V�%6cS%p������ч�BaNl"\��)p��4.L�٬��@��ʗ��O�zor҂��C�~��f#��_��p�j��^�jGQ�-Rh���C�R������U�댑/�J�mC���K�iI�Y���֥`�|���s��V�6C]@\=��T��F�$a�5�A�=FU�-I^����n�υ/'����Jq�9k�4B�^KƵ�a_��Ԉ����dI.�؅ �)���>m�����o_�7\y��F�� �i�_���^��e/V=����a�Ƽ��Гp!�WL
|��l�����p;�0�UՏ/m���bR:͟�ؠ����!ySהnǝ�������o�՝���Y6����7� AR��ʞ)ss���O��d#�˥N\����n�)����|K��
\cW(6�3tx��׈���͹��l|��;�Y����!:$�7#u��gM҇��;��*�ps�D���D:Z~T{���C��$��CW�羪����|H���3������Y��<�X����Ԕ��Uj:��G��{�х�����ø�
��K
���V[hE�b��
�!pE� �}(x��黜��e�D�����Я�&�\��W��)��"J^������d���}��dEY�v��rR�i�4xˏ#ib�<Q�F��0���0!��l	ռ�:�n�C����d�s�&��)R�K�1CE�=�[D�280i�kŦJiv-#����o��i���C���?�w$,{j'�e�M��>���[��������,�W��3X���ğ�e.H�޽��F�ɹn�*��Ș4/1)���8���ܤ�׿hFG�:Gu�W�b�n�ý��[5���
	�F5:S-��-�Mή5s�D�x��8�"�Szkm��..�R�O�P�Ip`����wkƭ�0��y��y�C�Fэ�#��3�MkҿЈ1�X����W6T}R��#5����t17x�@���L�+%x+V�vp��d]~��u�M�U%�]�T�y4ݏ
�a����.� Di?(�g1����z�ق
C���Z!˯(�WK�ϊ6�J:N��'�<�:_O�5�R��^A��3���W��0��-�WIT�s}��_2(�gR�3���
��$ۚ6��K�G�&q����WG����c�=/"Jjj��$]Q<A�L!���҈�������F��?_Dq0Q��C�>���?n7�e�Iȫu�~����2����_�1M����u�
%0��@��o�f�eJgB@�IuY�"�q�����O�]�װ��ݯ1H4i��u��ZKX>EX�˦���.?֥%�%~�h������]���8ȰJ�����:�(Dp߹kE��-���>;X��?G�W���ޱ�41���M�s.��j�zz���ŨM\�� t�F��z�u"�Fyr	��$���oA�9=��b�ԓ`W��2!�eD|T��"�n� 5H�9�,Qͽ�}���>سr�1�#�R�����I�<5cE�4.���"B���.ўL�s��@X��	���̠ζ�J=�k�������axű���Ǒ�R.߰F������4!�B����|�a�N�^�M���#e�Y�	�p���^?La��������h���l�A�Hb�1<��������j0<C�ꠓ8����ˋ�߇�3w��F��~J���<\���ǁ�{�����k���M�����~;nF_{��~Xb��jV)0:���$t�h,�K�"mӱ�����J{��� �z�)	!�͏M���]�y!w#mX@CF�_�A�}���Ϸ`�����+��l��ZJ���C�z���94�~��!�W0r����#�=z��2za
�
�3��?�5$B��t��Y %!^�%o� @�E7"V��r2���r:���;�_0Л.�1���*w'=���l�� ޼�қG5/U��g�/Sjt�s��`Y���E^��/�r>;�pwmC�UH	�z�<;�� }�Z��7�p�|ol�۳W����g�:%�����'}X@�m�o���E�9kE���R����9�/�
�AOE�W��g 1�R<��#v�p��9��1-�9�͖���"�>�r��Y��=�覂i��(�Y��a���L���wFz�r�E ��Ԛ��Hw,G�^j]1̵N��� ������G6Y��.8Q����@�� ��G������5|�1>�kIl*�#Ql�hG�D����qc������}��x�9�K,4�Wp���rG�����F)y��]1���Y�T�Jw�oa��p���̉:�1��S&��R��q{��ļ�����{,�*X�Q�?�������y����@7����$�?C&��Ǌ��(O$~~��� ���[m�)<ˣ���#נ��8��3���
�L��"H��$�P���_�u��������h��IT"M�g��n�y�
���!�Wx�����nu�WMƵ���g-���p����#qi��ǫmK�.XQ�Z�?聜<�`��t���D�и��s��e�<���O𫬈opӑ�:)_�Y�%ʢ�K�h\�d�*� ���z1#��Rqհ��p�ɠ�]@J3�$)�Z���x���=�m+�7����0Xx�t��@k�i��c*!�I}&%���
#Ճ�ˑ/��ת{��k��=�UT~3�}>Y�b��pA�� ��GX/BF䑊;��W(��V�����g��"��vy����/����1�����G�RSa�.�<�Y��z��\S����NA{�+� ������<^���P��JA�Q��)]���D=Fb�)4uy��zx��i�������[���h���M��\��0���I��I^#n2��'�Y�g�=x�_��e�yyG����XJv|���4��Ev�맟y��Kuab|�=�ZP�Vs{�V����lm�����(:���'u�4�/?F���W�r���� �X�C�-+� ɘ>�3ô��U�s�W���az��nܸa>�!�{U,ϩ�9O�
����@Z���J���Sk�z��XdB�lf�4e�+ۃ���Q����Xy\�TP^�V�%:����C��)���0n!k�S$����×�"3�O;����v3�7�Z�0ZۼvG�2�"�(��Z���;�a5�SxВ�s�~��Sr`���-?D�b�u��܉�wdU�/�8,C^�rN�r��G9;g͟Sk���&:\�v�>;˵���]�z�~�CGm�B��j
ԭ�W��ʧ�Y�=��y����k������f}ѪH���Fraي�"N�=HΤ��&��3s ��yW����˕����ot�:�9�-)۴G���b�/<�y��Y�]v�h�<-t�'�:�>���+𩁢:��#W�
x6�i~t�|w�\���Kk��pgke}�Ɨ�=�pZ��q�As#)�d,�d���C
w9_��AQg����ƫ��������O<g�Ѥ�N�]�+�nM�Q\�����r%E��|����Ǩ ��e����U��R����v��zZ*����>m>�G�j��a�(O6���Q�s�}7�0I��'�ݶې�°`�@ųXf�{������Ub!�kS�\Vu�G�8K$�OY
'9���s\�"=���o[�j��S�J��[)�������"��龒`l������K��C�����ڈ���BP���!��8�؋�nuy�Y;�(��2d|�n���$C,#�l	�M�┳i�zI��s�>R�V��֜_3^.=�of�8�P/��)�k� �R��̷��X(*�7�z�E�;i�7c��d���M
�2𜆈k,˫'Z�U& j��Nˋ�U�OPft���R{翑��%R4�*=XӮͷ��@��Dv�􁔢�z1�F�Yjg���&�ݓ���tr²�JG���=��l7�z^��z��y߇�)2�1��;zso���唛Lz���J׮|��9�V~�r�t+v3�1fm>p�$�\���u�qκQA�D�~�MN�qH�k�_g4!��������w������g�ciS�X?���_�fwQ��a���T���Zr��l��-J��7�Bu����|����S�)J����E��9����R�CÒJ�Ep�����T�'!Z>E���6�@[���q������O5E�op��ݪ�Y� ��
�Sy����3�w��d5%��/�5���o�(D��C�W�"�hFèc�f��&RH-60傑mh���)$���Yۗ
��cu5cEk_���
�8�p×^u�.uS�(�qF���nL�����"�wȋ%�Qr1������=��J�)�Ù����h�&��g�]�����{#�(�ې��	�<GM�[�E����z�/��}eb�G �_�h�2<���`؂C�2���$)��!L��lf5�U�]�Pi��	��ޜ^���P��f�r�&VFG�$����kc�T2 n���-�'[�$�F<EhoE3k#�.}�-1?W�({a+��a���\�c��W�!}#n���-_/$f�f��?�G�J$�K�G-ި�Y��6!��Tr�huR�no���kjJN������(���$ �����_e��$��뙱��D/Q��@4��L9��:�sP*zW$�"N`�Ԧ���x�L��u!��)�����#N�STn��aMb_*p$� ���;4�&6��g�V"i��j�bkVD���K��YE������%,߆�a�#�ѱ	#�p_M��t �w3��i��޿�9 }�
��i^�c�&��-l��VJ��I��t����P\���]r"������xe��o�4�P������?㩎:��y���͜mr3�s�̨�U�k%�y2h��i��w�"�����<�6�~Itw� ���GN]K��;^ ��Rm�>�dF���K|�����%����m�F��G*��/8���85xg�It��v�J��)85�{F�"�VR�%p1'OԸ��g����&���`��nO�A�D�
(���Z9�l�1w�{ �H��0�� �ݠ������½��F���}��J����k[��x�j� .)�*!qf����*�x	<W[广G���&�[��'%��+���q��qI�-w��iG�!�dv�o51�/M���h_���3v+՗�D'&�J*�&w��ms[�ǡA��"��]-��P
kz��mj���d���[��z�;i{ݝ⽇(�#ha�CX.1�s�; ��3���/O�V�����E�UNt��k�WR���U*i���b%n{$m�g��K0$�fm���My��,AcJ��IF<�;��0�IvVh�TBuV�4��v/Q��}�[��v���=��E�f@�n{�7�m V��-���0��@�i�C��H]p�у����W�/��.�����D3%�1~)�� �<ڦ�%���@���x��t��T*1�y}����Ow�)��k;7�Y�O�^��za�v���犆���7��??���d �9]E*@E����=b�	��A(Qh��JpJr}m�̞���^$�~��)��^c��<�!���F~5���p���1�$�Te��``e[C`h��ъ=>;�(§�E43�9��^�B'�xq+�x��6%'�����er�y�����[LxߙM7Fם�(�C*,�G����|�j�9|-mϑ¢��HZq3�Y���\@�|�&+
fu�D��>����.���e� �ѧ?����y�� ~�Og�ժV���;b��3�f;G��v9`��)�@�đX�J�DJ/�����(���$,�t����=��31o:�w��yWaQ��l������؜��5V���G������B�m�;��Al��ڋ���P�qP�m�Y�������r��F����^m�n����.v�U��n���g�Tt����K{��qr`��t���AL����2�؅�Z;��d�+6n5��u ��_j��6���h�/�v+e��5��2��7���ǷD���[�a�|�7�G�F�%��[v�'멲�nuo0¡�][��d����^*$xp
m��1*3�
�H9����rOgGl��Q�5���X�_֤v-to�3mJҥ<���<Y�����2�O�a=���Om�a���u�.7��y!C�*v5���v�d��[􈘰/Û>&x$r�D��U��-#���H�*�6`Rq��烈X1��^�\�b6&jBob��F�Ġ�Lg͌��S�j?��_��<	���ZI�!��#Թ/�\�N�4=���.�����!�ة��V�o�:��k5�l2��[{m��&��d
�W�h�=�&طtx�
_���#&??�$���!��P1��^��91?c(?a�{�ymO�b�E%���Q�y�I�N9Q�mf�$�`y�i|-Hc%ϑ���T�S'�G��NU�ZA��f��a]�1z��(�Ԁ�M��=*�l�R4��5ܺEO��_�Q�OK~\�V��5�N���桳����g��O~6X�W����B���	0�f�Eabm��'�� ��w�$�B�Ψޔg��|)��)�~l�@��ų�ݞͦ4��6&}�ͫzDf#A��t��^�A'�iMMaK��B>���lG�;�����v��7���ۗ^�~�-�딦��<=�ᾚ���U�`A�=�@�R�(������IЂ�Q��4t#ì���m��*%߾�����{����m�}�����Q�^��kI�֝���{��d�k�w�܍�)�p���bAF�I�� ����kT�F���΍��QSz�#C��u)��x�}[&���,ҿ_n�c�
�Y���PǤ��nK.���t���j�i�(���YYE$H�ﯮ5��H9�e���ǩ3��X-e�F!{T���Rt0��f��]��e2M����K�g��4��<�d]˽~�O�����7K�C��PDk�"q36������@�_�{7��W`PȟFg@�olM�>_��/�H���f��!�������ޛ��S�aHK���.�ܖ�Q���T��y��?�]�����7��[PN�ò�B����� �"c�;&��B8��bO��k���|�`l����/U��^Eu��}ʄ�8m�	��>"��sR1�_�	óEwf��W��!����5����B{Σ�/^�M�;Jc/���Ҧ݋�CT��$T�8��لZ�[B�ʺ���rt���(���y�!�y��f��z>G��̖E9�;��sX�$�a�;�]0��K0�ޤ��$��p}����]�=����&��9\\�1j�]�����4V�~����l��4C�y-+'��n����]�?�i��jh��Fk^��	��P��B�\��*�<�Lo�������b�{T�.I�%Ϝ�����S:�K}�L9�N�/~�d��	�'xT���[��zj4DD�X�	���ey���u
��(#ۅ�y���S��^�ч���x���z�WM���vh՟��~lt^*3�,�eo�2!~���'��GhZ��_�����6�R�ʉ��i��OZ�%���*��W�a*�c#�@.��_�<�<�כ���nAvL������]���l�d2��h��U��R�������]�g�8�Y�UP�V�����X���%I�����E��S?N%aK�ҠӀ����m/Y�u�<Q4e����tr�@pTX�PY�GT��Z��`�n>ܢ	�����&Cc>A��X۽�_#F�=��
,+��U��>��8#�3�vv��X��Wx�!c�mF=��sD�_+����F
a����	j�^�]��FFaT(QGBe�]3T�ʠC�dNg�B\7���M�s�*�LHu�y�;�e�t�����C�Z�(���9�8q��O���������Kr��:�:	u:C�l�c��mӣC����8
��v�s�$�-(�s�h�����d������ϳ�#��J�殉n�|����S���*|�����*�ࡼ3�]ͮ�rC�EY�P?H2�pu��a�����Js`�c�:�4N��K�Đm�2�[*7f���J�n�����t"+�M�Qb|��ư��)e�ϰ�-`��Mއ��"��^i>"c�1UN#�;^�tZб7d}��/w��h�q�����[fDM�B�0m&C (�mWY_$,��a$xA�ly�m�5xX��t}0|�rY���^m�������⪘��Az��s��h��77?�^��z�i�=�l=���\A
��Z-�|= m�3
���?�I�c�����IC�Ͱ�-4����E���5�Q]�]��R���R�����>T�g���2]����(?G (ֱO��<1��wr_����u�ܚ�����^X�2ʔ�789� ���ɿ�U<(�?13��9���Z�D�5���A;{d\�K��	mÂ��+6��#����s���v�]�-i3��k�V�zH)I�yg����K$w%�w�Z��o�_x~*fg���o��6���u>��v��S�a��y�o�6+�:������~v"9��zG�G��J/[�޹b&��3	S��x�zvjؽ(�2��m)�2�R� kT1Y���c?���ْJg�-�$��^DO��oH%"��꧙�yݲٮJL���}�r言���[ۋ�����[�z6ڛa`hy�)���ɑ9>�h��KE���\��tgi<��d��U�Q(�'���}��*��k�2_ ��\���{=}=�E�`.�2Mi�5���Ct�nq�Gbb��KɋS���y���Y@#����g������Qg��{`�~�����~�\lډQe�$�w�ܣ�(��]ϿTC��>�=A*ܴ�ǹ��fמ�hO���iTb1����WAT?B���gt#1�p��`Q�[��V�B���G(����atW�Yf��aB�\뚪=�����;B���ʁX����B
xҎQ�+Ȼ�,+#1�������M���W��K�MP������p̛�8a7{�G}-��e��7�� �3ן;�R��_sn��iɤ}y_8�$h8��$��Ru��9K�sa�jP�[��*@��iB�*�H��<��
S�CP/tR�a�ń�?�Ө8!�ju��:.e���_��;&�b]i�i[�i�����h�y��z��(1W!P�C�F�n�8])��l�E���������/3�&�$A�	�1)Ɲ�y�VF����WA�I��,��L��يJD�毡!4��큙f�S��?�o�� 8�9��s?�Py�X=���)�8tw��f5d�VO�F�A�~��
Sl"�أ�bx���ys�g�s�o&T<���F���>�����}C������*�.}o���q\_E��u��
Pt��0�[��'����~̘���-g���]6�X���C7�@i@�︆���Y�g�҇��Z���b�G!��kn�����/�Iҥ�\�l�-EN����2ɲL�gy+w�Az���\�2)�gWXza�m��Xۗ�+��M��[2�A�0k�Cs�� C*�/����^E�Xo���n���{����s7\7�~>���Yq�^ ؇":��~�/t�]B}�Gg;7g�k���n5�HtR�����uO���H�\��Q�ٞ?���2�A��W��BW���[d_�Ud:m��A��b�B���&K���.8�t�v�{�b�d2N��O�}*�����	��$����k/���t��^�����I���2�w?ѩi��ZXO���.��*�wԷڂv������ܘ�KM�?M� ��' _y�[ma�+_rTG�)I��?ޯ>������>�el��ͺ�9�P1�K&�J����`\)F/ "j�,ϸ���]�ھ/���W#\NQ��YeJ�P*(.%zn5{VG���<se٫/�+@1��`vf��ᑤ���):���A���s�W28���\q)�_��lڬ���{�����?P]��$~������Z�C���F���53���H=�2|�殴�qa�<�̐D�>ôoNa��V_(��o<6�R�رtwy�g�^����51��J��6l�T�\a�5g�����K�ћ����%j6�A����]�S�;���[�a�r=�e�yk�;Gx������)�/�@<���BT�F=JV޴9)�q�ꂣj�.C���465�N�~��{�}Py��&W%�ԁt�Fi��w5��Ao�*�59�����:ə{�,���Ő���P�K ��U�y��[>�3���39 S���kJ�ڷU��Y�Z����8N��o�����`Iػ�R���Üz���+�B'(^_G�Eo�Q(!��c)'+�8���7x�R��G��JF��<�ps��y�4���]]6��0��Ñ��)��1
�5�?$�g�Z�轭ء�3s����`U���10�W�B��D�O�1�@��H�u��;�R�1�tu���%f��:ҁ:��-^�#lQ�������Ic/�6�e��!���h���uv2+�N�ۋ�ad%�w���y�n��,���{AG������3�3I�/���n�I��Q����)p z籊���_�0ر��ٝ��"�%�vr�ꠚ� C?�^0���U3�)��x˰Fɏ�M#}y��#p��Z(rf���ݑ}#���<{���S�8�yw��u��x
�m�q4���ƛ-n����RՀ2���M�=F�S�lgmVCT���ߛ�9@]�����յ9�7�{˲����f�l���������¡�ퟅݎ�U�'(�w7t�S̠v��������+����*?��h�½;��o�&���=�� ��_ a='��Z�]��2�g�5<<=��p:��(�p
K��_�0�,��헱;�^��k��Y��� je!</�6�%�G����iك�N����{\����A}�����(a���Ə���φ�Q�T��1�ӆk+��Ae�f=�7n(߽��&p����'�x�������7��T����@�H�gkKvmu�ضhj6vIA?k�����_��FVmI�bt#�� GE�vy������6u�(+Ai���FO%���:��F�����#���-�+5�(+A닉o�
w�ID�~���w͊��^�L�K*�g��^����\p��ȶ,{"��^���X��8y�烂k)��й��� _׹z�Wf�3ul����'m�;{x���r+~�ܲ,������d���w�%7��^���G��+����{����/��6����N��h̨�[X�zu�ɑ��D��9>��\�x�Sv~��XV��z���Kdj���u*�IN�0d�3�j��U��|D����V����_��Y��Q򌢴a^�CX����TU6\����A��x��!�̆o@�����~��כ~%^[�o�"__o9k�D`*v�៺2����p u7��́nf�f[U*���D�&�]Zz�{ʪ���HR�j'����F�R�8kD��X���?4y�^QM�W��AE�WZ�)�9�p��R����[����z_ZeS�qE{�ŷN�J}�T^!`��(o�l>u�`ԋoGA�3X�,`�fg�4U5�!�)򒗄>Ӄۭ*|�cT(Ƕ>��@|ƞR�0�ާj?-�������>��W��f���ޮ'��"��nli@U��l8o�S
��"T���n���w(��kҰ�e%$._2X0^��ŗ��/�pIw˩K{@�rWp��30z>�`��w���9�[�������h߯1���ǭ`����2�Ɣ�ڐlS�򶭁ٟQ&V�]��G���n�3r%��tyE�8.��U��� ��yUϺ%���Q�+�⻹��U�� ����7�o�G	Y:��$�b<%7�7/�s ���Є��,%�&�s���)��%9�u�#O��o�ӎ/5�
L�w������{v'_@���*\�J]���6���p�|�4ۅP!"��wn`��=,k��z&ܷ�S�գ=����t���Ģ.��f!�E{�������-U�7�,��+���[X9\bZ��_{󗸝�%Ȧ�.Cc/�:�Y<�o��|	��R|	�z��Lo(?�﫟-L�Q��Q����N~V�x���"^��גr������ʣ{���e�r}3K������*��^�nO�;E��X�3�!#�&�h��̇%o_�	�!0�����X�K\�뺆�	���(K�FY⟣��ˬ�	~� ��N� s?��d]�,��U���jL*g8�1���t�z����<$��u6w�P-+�,�K��\�1V�G{
%�����U���w� �c�º[J����]�Oo�/8�����Cp���l��Ycl�~&�`s�!��xV�}g�/���s#��IC�ߝ�I�B�{x�B���uE��LV'��f��4��j� =���@��承��p�[��ط�溤H�����/�#���-k�I�[q�?!��gۮ��㈮�4��� ����1��{$�-��L	Z{��Tǎ�tH
t�u�E��x������w�0ؾ7�~p��ا�^��N�r+�g�?���$�kQ�\m��{����Q�����k�e
������Ҡ�:�kw�S��-��_i���Y�LĦ����7���e$�ύ���<��ب����J�Xr�WÎ������M��b�래睜����!�ԗ1Ihr���|ex�&�'+Aqf���!wɑTvnu�#�$�j�pg�02U�i�z(��X綩d��<�?���Hk`�U~�cU�uvjx<��0���c��s<�G!�e��S(�?N� ��>�v�fe6y������� /ГR�x��z�$b6�WI��g\�Dſ�h��5�c�g&E+tx��w���,o�Jj3�!1�5�����W�,~d^��-�1�V{��j����뇵3Կ�bY�V���=���̼�>�-�Լ-��R�!.��9�R%KǹNO�-��禼�;�y�Ч�;ū��#�u���}s_�$}�Bg�qj��~m�J�%��J������}�������9�����,��Բ�S�e����h���tq� �
u��.ժwZ�c^�~O�ҁ�G|��[�����õ:��6�;�e�K7
�
�f�?	(��!�l�B�b�����o���ޑ���p���؄ٯUT��Չf�H_)�{����f�,R�Qu�v3训�?յP�>���G��_,��������U�NA�����k<9k>���2����� ��K�˿K��d��:V�P^xX8��87���ء͖{��+����uzsW�����D��q��e�{둕��!�pJ1�d���9i�п4��c.����.q��\�����|ol���A�BgZ4�W�(W�g��XI�\=��@�T)�8���N�'�Й�[�W�w6S��܁�L��ЛЏ�J��s��'�G8��
��)ª�$�5�W.�N��<��sJ1��.�N�J܉�io�B���[�S��i�ſk�S�yq���;���q�+z��ii��~$�������v=;#h��Y��y+ �6}u�ɲ��C�3d�����A�n�����N=-ۭW2���u���f������=���s4��)��_���g��~�-q[��g��v�f|_�\�����JP� ��5���$��M�u�R�r��3?�qGG�y-=�H�0L0�?�p�(z%7| ��N����ܴ<M@>UDB��m�sQ{���'E~��3i��8���=t7A^ʨ8���
�qYm�p9c/�B����ۆX�(��L�8��8�ڷ_�)fĤ�/l�5s�y@�wH��B��$J])�ԛ)�X囵���'i�� �L&��33�K92�I��q���=��fT+���bc��O���W�w��%�4R�%-nW��n����軌����3+��k\n���uj|鸭�wrBi�_ެh�"w���.�oE&���s�]�!��=s6q��A���D�zCAK��`�2 ~s-�Ι9�5�P��)��Q�r�r�N^���� ����~��.��H�Z_2�@���7�4��L
��.y��{8�\3��57�!�3�ϗ���zHg[nn�$�Z/�6ԔG��k�G~^�|�;�l��7�3�� %�؋�-K��|um�v��
���e=����q��Dx��	$k~�����/���ʲ��*BL�����
�
vE�-(>�����|Y��i(��_@:��xv�$���"�C�����Wn�榊�����:s�e�̃�H�e7��^m��$ʿ;���Z����m_'1�@?b����#}8�������X��1���H���F�Ia�+,Sy��^��T��CC��w�o�/�E���-p"8Y�-��@����n|����0�a�w\k�WF��8yVH��m�� Ct^-j	�^Zd>����H<��<��m��WxL^��Q��3?�1"�_��1�_�56.�쉮s���	�@^��"X�*�K�f���N\)Ζ���y�)$NcS����c�	q����H�?n�Ϧo��|V�3X��p�m�]�n�d��́�����*ob���j�?�9U�)������0|cxO�f\t��&��Txq�����T�H�q���8�#>~�m��_)�G̽�����Fp��i�a֩�φY�s(����Ƿ:J	A��9�7A7Ӕ��R�����W`��3	F�@�RqZ�)a�k�:,?�����R*��|��N
1����R�����%��� ��{I�Y���1�[��Z��5]�c�c��kBj��7!�o������Υ���5�v���Oi��Y�� �D]N5<ZA�ʲ	@�R�Exʎ3�I:L˓�9Φ�l���ײ�~��.U����-��CG-<����}��qRһG=ݬE0�J�ν~��H�viI?�ֺ�;!�Ȩ*�
ߌ����(	��{��U���3/�O�0_dx� ��)���H"�!��y��/��VRF��S�Ђ}�����̏�wLwhD���V�H`Q�nsQ��g\�e��a�19l�UD���8� �s ɋ_������>�������_A��4�a�4�yî}�zm|���8}�����+Å�4a�>43���m�ɒ*���u��A���ϥh��.�{�6�	�>/u|N�:PN��0'@�7`�v>C��W���5�s��A�/#�Xm����"��(��gA{;|�kŜ��DeU�P3y���ء��0)�Q�Lt��������վ�4��8L}n�t��;$0#a��4ɨ�>3����>6��'u�'�U_ѣ�P+ŽlY7��s�F9X�y���Hj�]�u�`���ho��yJ�y�1�!�?�Qub4�35�u��($�sL{�"(���2-��&��|��1�u���z��"P�H/�0�� ���/��
ƣZ{���ӯJ��c�[�����IE)tA��D�ߊ\r���*���3�-�TnI����f��.�m�w��n66�����`�=o���yy���շk���S@�œ��_-ގk����W2�N��ҫ�ʘ�q��4�jݘ��S��YV���_$#Ӻ�<���7Jm��N��ʽ���	�ΘbC��M��®�t�<��\�	�+3��S��pl�[!1�0�J�d/��{�&?7(�>j���KߺZ��~��u��8�廇�,����\�������>,
��-����e�v��A�yM{����@��n��6.��8��읔�p�~��*^х5��}z��w��I�PO�vI|�K���2[��6�JN�jDq�����s>��^���"�{����)���57�
�J�>�4��a�Z/�A�pC��?{i��qԾeZ��tm��o��p��|�YLw��a=t#zp�	��\Z�A�-�8�� G=��wc�=&Y\���B/����g�6���*[+�B^�G��RmM�"Z��B�I 7�}�4~�#��>DR.�x�����t" ��`�0%�M�	#'�#��S��{m�M�k{M��mא L��j���K D~��A߲�P}������|>�y^f��_Ȅ����:������_,�
���2w��ʥ�8���F�Ӧ�$�72����
�q+��� s�����=��z�qN��Z��?7p���{d��+�9寍��	8��e��|�=�_uo&km�+qC�
�����H��}د���.iD4,��GZ=���}Sv�Y�mJ����c��)MSJ{�F���	k���ő0�О��o����n�{�V�����z�D�Ck����w�]cqЯ�nȸ"J�2͗4����f^��W���!�ow����M�L��r�E�A���nC�R-���Q���5���Ehl���웲��p8�/�X̞up	��
��DO_�fj��Ɇ�V`w����^�i���B��
�I:�i��|�9܈�nк5zT�G����V�Z�YbV�YT��~�������
ň��o�NWhmWj��z.WF}F�?vx�:q�[��S�t��U�.�@�9�tu|8w�6��� �����Y��QU�+WL5����S[;rj|�i8j#I�K.��%�&�zD��Q8	�[�>�<�K�H��a�2�˃�i�������p΀�t+pe"�c�DC���0=O���	� ��Vо��5���X?��ƪ���6.�d*�6:-�#�&fT���b(Uu��+�s+K����o��hس�nj@���c�K�D&蒬��K�v◕F�`��<U�Ul�)�������}�_Qkw ��3�X�֯�$���kH;�-G�T]���qw������	wx��0<�Nڭ�u��q-[�4�D�
�M���f�wv@�"T����3=!O��т�wid{x�¼��r����y��D[��Mj��6��>�/��0��t\�}��l�B��5a�c$O2��ގ�A4�k���]$�P[������ܯ�y�Y�-4v���<qg��,�g��D�4�=$����,
�}0ݯV��jޝ9��	ZOV#��Ӫ^�0;e=M^��jCk�)۠<>�������>xm�^���v�ab��Zϧ�*J(M-���<*
�^����Z���&pO�/Y'F�f�h�
	���(�ӯ�`�^��UMCg������]��(�6��s��߶��6��{�fU7�o��Õ^���z���@�����nf�`����Ik�E��n�*_��P� ]ŗ+%�dְƇ>O��u�����$���GE�ή� �غ��)�J�i�ܤ,�V�10�]�F�4����-�ѹ��+WM��-i ��H�ش��c�HD3��e�U��0>�0z��1۞����y��hq��S*��˧0#`��3����w��t��2����H�X
�z�<ӧ"�A\���\�����C�8����������vv|��r2<�>�X>D���
/"�q��X	��/�~7b��	�֫�a��ղ���N�����y˵��aF�u-u�z�"&z�Q�B��`����M���F;x��P�	%,���S>���p��JE�>W�}�t��X�T���ɿ	,Ê��Q�}ءj��L"U[�s�e3��Q�o7ܹ'cK��͋_���.�e*)�_��yB@2I� Q�P��<O�)���7#�bw�p���\F�<��3+�g�GR�,,�<�[
e7�薆,��xu�ŭ��y��U阖�>�@۝粉f�����g�˟���Lh
�u�=0�O:h~��Ω�Y��;�R�eK|�*�h�lm�kA�у�����,�&�?���|Y���/2��&k�Q$U%��93Hi
����Nl[Lgܴ�^�)�� �&f�����$�YfrE��M|�!��(�LK�p�t�F�)�JG=���M�'�M���U���p+��V�qݼ9��ç�Q�~�3
��Us��6�t��o������*f�� ��Ӡ;�ڡ����n Ng}�0�H��Zyz����Hw��E=?l�T����Sl,^#�+4��I�����$���y�c)\%L0�k�a͵a�d$�4bIiq�jЖs�0h�������r�u��}3�*�ګp[��8i�a���F�2uRU�m@���&�8��Ec���(��n�j9�E"s��N��q�d�:�-��lx���ψ{�L8�~|�lCمnǸ7+��0ّ�y3�I�}�T����ދ+��?����?����(��Z�"t��vt�+�m\t��#y�����?lR�o�@C`�ݮ:bv�� ��Pd'��~������1���	�yk����r�/̂vɜ��Z>$��lt�u��1c�!�t��eVU��#�t+<��ECXbc����h|%��	l��ô/ ��?�|��-�<u%��u1<�����wc`��[�*�ps�4���SzK"9�E>r�K�Qb���\k���
�㘰w��`.���sY�hֳhi��VM�.���Eq1*<���ƨ�I3>���w� Jv<���u�z�߅}��$55���%�Q�I���	
P�f�w3�����g�l�ߙq͊~J�{5��71p���ZR��4�Jdb<,�0ۦ��r�!t����Sf�� 	����-���;fK�Y�7���n��9Pf5�p~��U��Qowtߏ�����h�ߨ�ƧR+U0���h1I͙3qq�E�=�׫%�A�ּҲ�fS�#�(�~�f�<��h�V\�8�F^�b�:�r�P��f�$N:�y򷞵e6z˦�<C�f�D�h�Yt4�%��`;��&3���Ο܏)�����"m�|�3:�r�w559e
6�Jճb�i����9<�\�����v�j~Fh:?\]d,�.��#Z���ּJ�r�c?�`�¶���ƍn[�����`���G&��	sg%�������V:����s3fuЂ��"��q�F6eBCi�і5̈=�>$E��ne0�]4*�$��t��Z�T�c��yܱ-����J/^&u=�p=��p����!��e�,����Hm��+c�58�J�寤�bA���!J�9�Ѩ�\�M!�Z[���'���>�@b�cu��sZ'��{� H�~���۽�<��V9uR�ɲp���чHJNS�#d�N�b&�p�T�P��l�\��!��\�F�n��8t0lڻ�$i^����]^卌����C���3�2CcMA1������xI_�?2O9']
p?������p5��V|4�W�ݝ�1�n�Iw�:���}9L�����
�-t� ��~�ͅ���ͬ�0+)�ܴb�}9�sV�;��۬O4��&$X�F[ƛ�T��.��1y������Af?��N+"�I��~S�Q6N�M����F��]��R� WKğ�Yi�҈/\n�P�=�D㚊��En<ڭkfL�nE>t � ����3�Ϩ�w�,kY�V�?��̙�.���Gy�p�M�u�t�7JH�!�#���g���'�%����y�ױ��ԫ���>q1̇�B �Abu$�+S'�{�L�N��W	���Z���]��LqC��y�x���*�vw]`�m
u���3�G0�
�$�~���W��}�y�g.�����2ieJ�g[�;�B5k�dk?�������^~����4�Gm�R��p���:e�J�L�+�y����z�ʟ���9'��xA��=�͇g�� T��ڽ&�(B�hàF׀t^-�o(�Q7{M�3!����tw�`׀b>~�����B0�9Кw��i׶��P�掀HzP1?�-��ea�W筮u3M���)�׃�A:�W�g���<^~Jq��I�%�q%�]�� �~TN�F�*�T���vso�E��:�=�@�1U}�EO��N��gR�E�	��&R������Z�ax5��$&ihb����{�	��SCUs���?�ǽy��W��f�u�oh��g�xG f��@����TAc���YpL�GD,�ڮ�B�J ��W�2�+�#���=L�ιY	㪔^S�?�A�x���6xp�M�����
����YoKL戇�-�o`�97i��4��x4�	O��߹Z����v&M��"k -�#�CӨ{KR70o,�)�����es_�N�x"ǼN�/5��֕aXTb���ZN��
���qr��o�d�9���y�e���'d��1v=�]"*�A^R,�~h�Ra麗�!��(޽i���G������k<v�@�Q�t*�uu�L����#����̟/�v�Z��a�pp�8��S��C� �*�c{�����
z�U���u��Qa��]� ��� �v�n	W�1��9 ��h��4RZ�G�9_�9�_ɱG~�IH�.%n�)��qb`j���޻kZF4���<��t��,<��F�$��:8hz&ϚV���N��GvaGlA�m��$���9����̒ݲA��}�fE�����Ē���CS�=�P8w�%o�X �i����/I�Z8���z7T�H�u�	u/U����U&��b$]>��l���Ks�/���K���1�_bmhy�<-O��>2f�����i������A���eʯ�⡢Z�TRx�2��������V��M/$��vCPe���:d�2bO�vu$���z~�<q�W~]�:6���9�&��ӳ��=�22�)�>�ao'=��}W�%���:5�����t��.����^n�z�J�cM�Ug>��5��.<7�n��MW�p�@OP~�+�*ީ6>0���x}�R����/��X��Ya!$p'ҰŊ��ЮI��\�Q���
�K%2.��=-4]p��h�ZyRM������ｖ�A��<�#�ppYc�=�I�S�	�֮Pq1�W9�k�v����U�`v��!L۪҃��4e� �C֖=�15���k��#\��R��dP gt�w�N������͆�Ǘ's�;���e��3`<�jl*@��xd2��Pa�6l���6�>w7����;ƨK�o�R�fp�5��^�%U�̟'q����Ȃ^�����b/(+j�)n=4��V�e���(�����9�Zzz ���:.�#"ݜ����u�̿���U�.K�!��
N�D�������WD$�
d݀��V�>e_�Т˦%a�f�p�a����9���'��y�]fKLn?��|������"8V���|O����T�7CN�U��ݑY��4�.�y&}COM,|MJ��ּ���tG��R=d��D�nʰ�/k����=@�f����M���"��ϰ=nW���_�Y"����W�!h����ݳ���2O��v�ԛ\>Ԩ�kJ��1�����b��egr���w�Ŝ~�f��+i���u�c��5)o��H��U��Ž�$���P�-8�[����+V:OW�]!�/ĻZj)$�_�W����#dH-%�m_
p#/˧����Z�<��T]�\tc&���E �*� ��p���$v�'7Z?|���e�[�n\<� G��T��7Z5%3�Ft+�i%O�?7�[2��;�%�����5�ݻ�ء��K����
��g�*��j�ۖ������Al�%'����BA�ڮ�n��G��1�����_i�+2�nŸ�@s�����I����o�'����J�*�)�o�=&���)�H����Dy�[�.��z�r�v8Li�`QC�FZ-N�2
V��:��mЪ��B���uY�
�NN���HM�D+�]=��ſ��	g�>�|���]/�fѽHW���CevҲҷ~�I5Y5�ý�.�& ZEi�[q�ev�wR����WG�h��b"33���{�t��
��i
������M>��/�Xqfl�\VI~��lm唸���,N�bg��v�,��f��-m�;`A���d��k�9پ7�م�V��Q9P��d\]�9��]���K>=��W��V�ꖷ�Dɠ��1��rB񺠾�U��[>���P�_������<�#	��Y���,�y�;�B��bψ\����c�R��Y��R�Je�LW3�y�1⢭I+�����Ւ97+��)jjE����jo�c1�%�e��gN���޷*=��w�@�'�T�d��Mb(暴�N�}��>��k�]�r�ԋ@~&xD�G�N%O9es.�M�.�ie��Q�jj��nc�0bo5�k�{��V�hgԮg6�{w�FD���WQ69�x��U5����+��T���/���a���30��^^`A$:��aʃ�8��%�����a ��ڗV}�8�-_H��s8�j��!q7�6�"8�-).��ܭ4�q�w��;lH�`�w�Re��������o�!6P��%V [�����-Z\���v�bg�p�+܌&;����xH��A�%�G�E�ŢS;�*��]N�&I^߭	N$�5b�F�>�@�����w�������~������%'��ܐ~�!�徚G�W�soŔ$�G����g#�%2�]�%�Q��D��[����n<�ޘk����
�r�
)��ؑ�jw�y�T�m�|�J��G�J�_ǋ�z� 1u����(��C�mY�t������A����2�䗒_��?�����P��k�֓�i�����eg QC��\gB>,��/�Bi2�~��#�Z����߃��;� �����1+��|�E�!���l��[y�t�Ή���&����U'E\",2�k��)5h�0�]���1��S�K��Z��Bk�z�F�T�y!C��&7���k^@�l�5w�.T�m�Ò��t<qj����_�'�=T%���@�uå"��N��Du##�6p�q�{6Ӕ]�Aف�]V����~P��1g�0!Lk���4�󀒣���:v����YV����q���d��")8�/ ^�w}��U"T�T�$�w��T��[�5r��B _��sQΤMz�:�Z����S�K�P쯇��3K��ۅ����K6��l�fkGA�?lZ�b�r�v s�]2�߁ϔ�����U��c0 /q%�cDu�����`�J��*��"-�������]wG��<�{�� �>�n�ާ&{#������{k�G�Wz��S����U�SS·Z�.���i�:HQ���L^
V�R������7���{j�ΈF=2�Dᙎ#.�Qd��;t�]Yh�p)������=�"_��
`���:����wW]��A%[�bO�^n�"	l4�s�\ٳ�^te{���z~x����"9#I��Y"<��	��jZ�)ů�B\��L�l� ��y���^Ƿ�1&���_b�;���)�^>��(��\D=»M����	6���q�@��c��)�����/�Ctk�b��#b��i����'���'���s�b�d3Y��K��@��37<��������%v�9��xO��{�Y�_3�k7GT!�ǀ��;��kj�J�1�r�G�_/��qy~x���DkL�X$�ù*c�,*����q�����C��yr��/=h��z55��6��%'C�/��)��Y�K��0�ܼU,��P��ʙ�� Q��V!e�ba}1�h-�w�����r��#"�R;/x�����]	�\{9d?BϚwM�0��2���[-�0牨�a��\}����m�0����T^9��}��+�t�꺶=��7y��N�s��e+� T&�د�駸B|�}��I��s����{��ꢠ�ּ�(>�˂�QS���TYh2s�g�nݿHg�#o��l�C�Kr۷Uxc���S<^xj�LT3�T)��*{��y�DZW���/&�mT���N����p��ڞ��>�Ľ3��hȂQ�(3!��c�|�!ǜ��	�1�|����m��,��Ϙ��zL�t�-��ɚ��"+�*D�c�����3�(N�d(�����v�����T3�\=���k5����O������Ԏ���}�F����t���w�*owTݧ�N�jϷ�R�?3k!�T�C�mb)v1�/�Ű�}�zZ�����S��oт�����b�-���C�� �m��>J��O��Hr}��R�R7�,����)8*����F;TMc�B�BUb�TkiA,���Ѷ�7��|�;W(�T�|ܲ5QI����B�����l��4��G~��W,Nq�0�$Ta��Q��%����T����m�+3��G�q�z�>�$$���(���F��A�%ڐz�I������<�5_��ִo=r�޶��,��?���V��_�0���l�h~+�F�Խu����wN6QOk�<��<qN����ep���åMf��*GI�6+-�u��"�k�D�{�$�\����=�ygC��Z�^�����d���<�1������w!��9ݪ� �3��;��ʽ��<� �-�O�?7w�Y:�o���?%�_�<M��S�Q�6�dT��Eo蒮�5WD�\C���455*x&��ZĚ_t��H�x�:,)��,�r{��z��h���oΊng~�Q����*﷪X��T�GP4��Yk�\b����Sʪ�a�7�����t�6��rϛ[�mJԺ��4�)��"723!O�����ˮ��=Z�E��|q�*�������������V��I�cH�嵽x~;!g��#��{7���M��#���R���ǖ�l�nb�� Ή���݅��.X��8f*a`*��
�wC�� ������aI�JK1�{,~��W;�wq:W��w�L���'�k�'oB�ӑO>3�3M!����M隇m�a�Y�l�ݤϋ�58��O�77���U��?Y�9t?3»�8F��
2զ��h�?��F�{�?��(���ޚD�l[j�L�ÉٗO�>�dm~<x�vk�[l�"�+(�"CwG�t<�X�Nh>,L:X���v�C�%�浪ϋ��\�������N_ ��ٜ35�����j�/p�^h�m��{d(�I�L!���L?+P;�Ny�;����RB�(��~{b�3���a�x|�����o�s�ܮE���r��)?���rI��Ka)G�ւEC�5�vZN�������#G&��g�n2n��{e2�g�<k���n�Xxκ�I\��A*8��W)-�"���Ec��*��ؿ�UuѪ�Dm.Zl���Y0�W�S[�"�dq/YS�r�4���J�/{��#QW�w[����@U���Q~?����j�9�}�'�3!�r#�eء������m�ҽ�X+׳��e�m?��Af�SfW���G�c�j�g�qH
��_��Jl�3�Ü{�k�k�R�(P_Ff� �5nټ?�VL��+|!�}"��jbO����]������o�W�u��Y��c��o�
1U���H=�/���}Q�w�zԓXv7��=%�d�Z��k\s&�l�=��vô=�Q���Jq@���;��K���y�/.����J.�'��~n�οiW��<%e���f�X�>�T�(Z~?��L�Cֳ7P��xҳ�x9v��W5��x�8_�#�W����p��Ibk������~ďęb.�dT�v�k�S�Lm�z��f��@`_��l��e�����jTL����;b�rt��cuxke���o�{���c����V��`��~���$ϷU!	��d��q�jdGJه=.@JJz6vܡy�����[-������}���w;;�ب@����WZ"3t�2�]	_�k�	�q���Au�u������(ʤ�ۡU�N���ve������gfS��T����;�4�'ǂ4���^�����r�?Ƹ���4`��c�%{$���EY-:�����9�SS��2鼝����(C�6Ky���>�^��'�u*lRb��$'�ePe|[,r�L���(+*q�X���2�.�Z"��p���T,&�J~;^���H�*�|5�Ǧ�2>Őn�Cͻ�C�HW��R8���԰�y�g*���>���FJ�M��Hjac�(�]f�V�K�dٖ|Gm@h�~��ge��GC�0k�m�PV��u9�rQ<��JA���@�[f�B��'TaN�p'�uԳ�,_��"yE��0�	�x��y:�C��������LWDZ�?I�:,��S�����]�����k+)��:��$����L��儶�82Gfx�A�[OzT{�|Y'a��M",�<�[Sfz� �ij0:��ͫ;H�sAV�G�H�p�!&���J-�z<��M�����xn`bpKqe7���k�ZR?��g����K_{(�������:ɾYM����Թ�v�D�5n��]a��u_�C���ez��g����#���(h������+93Q�q�Π�I�{ʐ5���G���o��p���2n5����O���P���pqC�z��h����~9��t29T�-��a�]��+{���a�����F�_��Ϭ}^�@��'}}�;��Q5�n{eeY��x��2.������E�*Q�}&n��Ģp�����u�<�_���#��w�R��'���n�\���^�N7]��D<�����������g���A��Y����_�W��2Ng����^[�i�<���/t�E��`|3��U����Ծ~e���=�������Ji�M]tJ�Sիq�č?[��\2��?�S���0�F�d���-��j�B�!��Bē����Ja%u���0x$��0����EB����w��K��'_{x�j�<N>ξz<��nW!�ٻLt$w6��)�h���y�#�(^i� SsCJ�EcE��|iJ��Y��9�S��݉��[~�_K����ez��%F�C�\v׿~XB��ڂ�?n��rI�C��[]-{!
W���5A8�,�gN�$��� �S��	�#���JZ��B=:`{�d�f%�(�ʬNac�j[�S�-��M����-�����Ű��ѫl3=��i����KŪ7�.!.������y��}�~6��&�n�ϱ �V%�X�{�����du��#��>�����7���?NG@���/��SK�"�2Cϓt`��޵�u'�C��F��sth�g�p�%>���2S/x{9��o�H�BI��1����h�vW�n5sx���E:��⹺�F�]��G�����ȸ��Kk�V��"���&[�S{DHm�PG�!�#^�bǑo�3詳�
���V�<�~$G�ߖl�o�w=������B���) ����|�m����L?�Kg�M��p��!����N�1���}�����FM�L�X�L�*a5ȇj�C���ԕ����4
�<U	䌂h-�Zo��.�xJ�{�����E�1��k�3��$�r����>��V*pOK��?� ��,�>dg%M�����pO�:�!�\�ӻ�$g3�,B�vӗ����ͺ�4�wV�G}%��[����08����&��zS�-��%
߹"�g-���p5�V�f�$J�~�hc��Ƽ���[�8����oK]�Bpi8��e_��־�?/�	2w>1?��%\$U������㋕����Y��y�]���T/qr�PD{�^�K��#�0�K��$�il(}lZ�v��þ�=3t�?��2���vj:��F�ǽ�D2ޭV�PP@o��6�	]iy�����!�xL,��E�Ae�? O���c��Ik���:��)�	K�hg	�8��e��oM�7�_RP�cp�����OK��D��5���m�W�B��KAU�~�L�K���Sm�&V���%K���]�'����4�u!`���s�Ç�7��0�Ŭ_�k�8o��d�����s�%���Fr+��K2j��
�*=�RD�qLkͬ�.���8e��U�b�%�G��{�;�O9l��EN�9�i�O��*Tc��4W� �V�}�Uތ�2�T���cp)!�(�W�ֆ�m��k-�����}��0Wt'
�#���_��bJ���~���KO�nr����qE!�~���3��e�ɟT�����I?5��8��{�;ߤ�]��s�ed�b��4�r�RZ{�fa��)���N�ZJ��^���ڏ��L�AG��	�x��+~ �y�;�5q�����
�-���m^�qG�7l_%OB�V	C�L�GQe����5VZu���jȑ�U��_��>��'\�al��^�h��<�2��,*3�u%~���N/��U�Gu�͎���˰rDK�>��c-�y�˻�FE�
��p���������L���,K�ݬ�O[%�3i P�ɀ�+�?��2.:Q���T���A\��$�_���-�V��o�p q��%[�|��ԛ�����B��sF[= �X�8S̤��ñ���E����ߝ�4~ᅝ��&�O+��i��ݜc�<��c-�Zh�/�aW^l'��F�nT|���Z􋿩F߾�wP��;%���N��� W&B�Q��A
�dd3�v��Ab�:�6�X>ޓ�$T"�(ì����B0������+�}�\=�%2����N��|��Q�SbкK&vR�s:K�w9�O��c��C����%�$���*등U��ٸAzI�̟����r�D�#_��À�`�aQi37���������al�e�'����>��� �T�ব���l.���3唝�>k����M���ﭭs]�X�w�6m��F���/��f�$M���=�2�&#*T��!�>���)l
Ye�?Gn+��!w��u?{r�luC��uٹ����f�4�譬��f����`�0q*^R��z���M}�lݾk�����m�:j��q|=��)va�&�]ԃ-W�����0v�y3�B�Tw�<�fb�t�M��`WCLZ �~(B�ޖsU���έ�a@s#+��ڢ#m�&2�H�zK#=����~厘2����L����YYK�@Q��:�uuؓ{%?�����Z����/�YJ<���R��n���u#8��'Sf7{�5�\ʵe�~xc�'z���y<x���B�'�m�p�:?]�ws�V�����n�\v����^�k�����l׬�'�?*fi'^�G�xP9�I�Tp�5�"L�G�o�t�s8w�m;��5��1fUy��bu��$��$�~��P�C�|��\`�e���B�g��K`g_��@Cb��c���x�׆��Y��W������.��J�.W-|�njPrL��H:t�2!u�A��#������[�6)�wm���O7�Z�z���ˋ�s؄����PK�@�M]�<,����u�p�z�p�V�>@��B*;'�����ǃ�i-���OEfj�EYF�x�[<�p�Vn-ss/D�L�(	@+Ty9 _K�*�|l��ِē�}�hF$�̥���v�z^��j(�(��qc�r���uU	a�y����o�����JDӆ"n�^���#e�z�Š+����OT>��U����GIu��`H(�Z^=��ВH�,8 $}D���á[w�����4�Z�&&��w&T�aַO�.L��y�#������i���X�sd�~�9<�[g����2mQ��yP+��5Th��߀��s���ӻS)�r��En������
��q��OH�(<��Ow��m���	��H�uSJ�~ݨ8��2OAd�$�/�Z#ok0�n�\g�8|o�����7=����u�M�	`�}ӹZ+%y[��Hlwu�`�,��"�.�&���[����?�ܵ8XWOY��L<W7e
���{8���M)�Y�
���}�XÏ�o�z�0�(�3�ڟ��ѳ��J���oh���~��z�����������}9��z�T�{'|�dPj�0U3�MB?C�6X���l5�H�zrP���] B��6�L�=Q�h�pF�/��b���p7�&8�H�-,��Vu�������4��֫����|�šM�?L�GBE����0�p����K�����P�DT���إcZ��R4���[��F���eTi*���d�5"�:S4����S|S�!�և�[�?�2wy�)ōJ���=δ�Tg��V��g}<۾��յ���SPD�����#��L�z1��m��v�a�|UP�g3ZpOړ(��;{�C�[̪r�â'O���pY��ZtFFG=�?��A@��q�I �.�xX��~ֿ��o�%��44;�*a�>�w ��N#m৿�B��]hk����O_�8�ktB���|ٔs��,�����Z� ^�� m�D��Kho/X����^P�"q��L�L^��;PO��n��tG���7�y-C�-�7W�
ݨ�	r���m�6U�H~a\���ݯ�ه���w#o�Xe�cN��ޥ���<i7�Ӹ�q��t����̣�I_Ğ�{��^�����ˊƖ�.�|C]M�ޓC�	��F�����z��ҡ'�F���UQ�7����ޕ�R��Qj/&WD�9Z��`|�=Ҧ�o�O�h��B��UZ.>x_��}��}�a�y�
Ӈ�<a����O�Lb��%oǐԈ�2��0\
�B�r�g��K�9X��<��l��`Vw�{��`��تm$�E�+%��b��T����T�c��	Y��*؟#��ْ�?ޗz5
��ϛηu��lߵ���p���S�R��h����~��� �5� �΁�O�]����CY�m��x��8�C�8��f��\.��"tJ���g�A�\��F���z�$=�4ie�~�MNN�+jD,��f�s�,�����Ĳ��bj��^ޝQ_$?³ k���IS�N���DE�x��.�6
T^RtuOQ%*Z%G��\�+��Pq�i�"G���d��.^��[^�˖+XQD�uJ7�Gb��lFV���t&���nxi+��۹����0KR��a��J����~��7�m�*d�ѥ��G�~�	��W0B�XoN=��iS���Wn�x�����{�Զzc�d�gI�՝��U����FP O,��һ���F<�c��J|�_"8(���YY����I�`����]�"�1R
Ҧ�P�@�k���<n��S�M�:�fyc�hT�ͪ��y4^+[��,y�ȯ3XgzH8�3Uf+p�z�kR�2L��I�|��M@ȟ,O�gĺ�����Ĉ���j�;��=,eF������XB��rb�h��Ƒ��s�a���ý2�޼���e���t�k���s=i���9T��� M3�n�\Y�^�]d��l ߍ��B�srθag��h.0�n��lwV�_���%�r�vuK���z�`r�����s�ME'�����Z"k��ʂ����Dݖ.�+t8)btiR�C�턗�hUXi�~�3=�j���o=���F!j�����ۇ�u����P��_y� E��H7��f��z�9��-�2�I�:�Fw!�`�3v� �_q#�`?�/��f��X��V�Das�3u�d��J�'M�Z���DJ�����z� s��En��z��1�}���pQ���C@������-f�
�4�}bϿ�X�VYM%������P��7�b�����w�-���i֫��Ul~Cح���kPL0<\��p�'���V�XA��3'q��k$���밚��S�%����������m-�6�~�C����C׺z�+VF�6:����q2TN�y�o˚u���>���u�"���E(�(�;��m�M�-�l-N�욇�;Q�ݶ���N��8חp��P��3��Q�A�ߴ`����݉�ղ�i'�y�]����>�l�T���D�2�VUʊ�:�?+A8������_����l��ʥ��oJ���a��'8O�J6��pwN� �dŃ(��˸�\�������
�Zq�z�.s4��ab42Tփa���c�.�9h�ٝ,�I\'	��^=a�2���~�"-N�P=ӗww�}�[#d��*x�ɅZhSVl6cS�U��*q��(�� ��� ���g�/
�DAG�#�w6IϷ���
c~�{fv�ߏ\"!�=!U{�W��v���jQE}��V�(�#� ؠ�8�l�q�����R\/�.1`Zbt(��D2��[��3O����/�|�e���i�*�����d�ӏ���A*��W���f�>J�Ӣ�	�_n�퐳7@O!3�]eD=� I����#��'q��efQ-�ט���J2�I[F�Ν�����u�c#k��<}|��kx�c&@���;� (�nZq��#����^��Ѻ{�v���=A��ΪX�4z��]��̮�{��Ɋ꫒�S+}�F�t�Fkbϼ�E׈(�t�@*�Z�����>�Q:�[���^���y"~��cJ����=��S_����ݮ$*		�B�˾�l#kBd���-{�${e��d��"{vc����1v�S�������s�u��:�=������X�C��C�U�@�Ild���� �t�D�R��S��Q�\�τЌ�Sl4x��N}���9U������_ڹ%R�!��~�a ��?�믬#�6'�oL��
*!�=��w~���k~ZS&zc�!Y뜗������a�&?$��G�ͭE���a�,���
A5�"�Ж˵~w�h����׬gx0}�J������ݭ)+?o�TA)�q��U��}p����A�4F�������`�=R]�te�4��R�]r䴁��y峥���U$5E95�n1f�[e�El�?֫���д)g}�͖�}g�'b�W`��K�З�b!��43JR5H�۱��
��q5�8t�TC�+q8�`�eQY�[�:&)�9P2]�X��<t 5w��ƿ�s/��f��)��;�5�n�h��t @���mȩ]�Ɲ6
�m��i�>y|�(rJ���u�I�d\:v�r���Yv�x�vYG���«�
��] ^?�Y�u����]F��v_>�(z5�Y��ݲ�-N�y�fh௛����,��e���\k�@�!{@ۓ� ��u��I������]���a7�VE��@�"��Id٧	�s��Va���K�bz H���mߥѨ�?��Y6�{z�;���0[s��� 6Z��Z���21�y��B���iV�e"� Ǩo��������]�Ыs�bu"�ܿ
J�^�� �04g���7v_k�#m�̦��k��ig1(Ԉ��i��NI.n��d�/f]�ܟ� 9g�eCt>�x��!墿��kX��m��&AE�9T�BW�D��HF)����f�x�{�hzNo�k{ a��0o�Z�(ʵͳ��a�8q)�l^�J�3-���[�,AkLf�s�o����Ķ��v�B�i�qg?�����$%*ϑ���%��HF����t��	)��Eco�b��.�K%E�c�|d7#����l;N������\\@�_���惽|?;��f�����0�R��-�|g����\fnxxʠ�2��pJY��1��ƙ�H��P��w�++@��%1���uS~����Z3Ɩ0D_ӓZEy̡�x�޾��(�}4̋�3M%�%#�6�왷6��ҘS�
/� ��,���� ��!�D���U8=W0eNDz
��~��ZG�b���/�р	k�Ը���W���'/_�Ř�y � ��:��*S����d4�+!���,{6�/�:x�-����<R�����Ա{:�p@�3U�c_���/r��O�D�q����#��F��;��x8���q-V?�j�"Y�.l!{7�B׍(.�,O|����ǎ���i55g�J�Ƒi��-
Y`B�+9���#��T{�8��� ��/�^�p�- ܞ<\)u,/�;ݙ�L5����??�y�<�Pɻ�|IC���B4����&WZ�D@_���Hٓ2�B2L-�h������N�u]ij
��)&{y��4���Z?/��y��t*ʸ3�yܗ�k5���v����� 4�h��3��o_d�QgL��n�ݰ2HZ��B{fn���Z5�VE�Hq��3 m��
O��mЗ�W��)Fu�5�����`�� .�/z�Ӂ��Ys譺*F��v6��H���g$"f����RI����(K�OΌݨu�]�����j�
��;��\����F�	�k���J� t��kP�u��ñ�Y);�@�'��J�G���Mo�v�z�~3��-׵g�}9���)��3],��ވ���@F*~C�ʏ���2n��9�n@;z�� ��A6+�۳'j�X�\�&�:x�Zpc!��FOP B�x1Z�ؔ�%S�"�7���wb�ˁ�$��ߏ����/�\����[�{�.�\�,f#�K.���w��B`3�����	s�����W�*�E`�ޜeϪɆK�f�F{�B��/H�w�&�<�n�o�<Y�9�~tT9	�5�)=b|���ߠ��w�H�Id���e}-����|���0[qΕ�֡���t ��J���$ꏕ]U�?��	�Ʉc��)y�ys�T��eo�B� �{�'c��:��Em��^
�M��S�-v��a���v�ǝׂ�}��n�aа���=<���I��npf�Ǒ?t[(���6�Q@��9�XC��-�R3�����g�r;����Vv~��"^�wcfm�S�X?)Nf�]r6�ҞLk��l���hbto:/eYZ�9�r`��זP%WXX�#Ɩ�F'Nh��ٝ��G{�A�j�c��_�͟�&��w�Vo�C���a}���N������"�#�ձgSvZr>À���U]ʽ�ï;�fǗJd��8#��'�ƿ����Ӹc'��8*���a�(����k]0iJD��@F�w˷�ձ݁O��+3�c{P���U0�4��J�B�R�j��A��.��p���E�}5 �Ž-�K�΁���;��&͔��Ə;2]���E%������a	{p"��r�	��-[c�o�o�ىI;e�ٕX�խE�l�>'�����Yr#�fA1�UU���pZ~�3 ��.��-�	��m T����g�P)�݀��i�1�_I-)T*����(�ߐ�f�wj}���	)�0�G��hC��/�C�����vt���C6�F5<�PĞ��?v��3�y;�⼕<
��R���g2̒�<Bn��H�=�X/�2{��TK�98ٔe��W
NN-G9^����ϟ�ZV;���(e-�~��J�+�t0�t�ӛ�Pr��n`&�Yc.�ҽ���QE�3���ˏ2;b�W�1`���&��<?��tx�y70)հ������N�,����lb̻ZK���ՠ\,:�9	9��pPD�i�c3��2��jM��##����ٰ����U�C�n|�ErWS�ٶ�����j���4�+:y R���'��lCK",��\?���mg�'l��3a�ЬXhK��q�5��f4��I�m�����p��7"OzW�Oy��>�-%�uc�{�E�t%ҏU�k�I�=	�sŝ�?>HT{�
�o��\��2���F��[YZ�Y�N�8S�7o���`�~|���8ǸNV?�oXz�WK�� ?�R_Hp��Ċ��3�JԂ+�Q��ڻ��}�������#�9t�X7���<��W7fn8|�3p��f>(t���
��9��?M�O�����6ۡ�FO�$�-w�C��(~5叹r����C�Բ��ٖ��0��V�!c�5Ln9�ь�&~��E�K���9�KP��Wϫ�±�03�:\գ���8l�R*UpUG�0s<��|
��v%�D�;���!D�R���[&���E?h�[\��?�yS��˭�Be��1�n��A���H٫F�4�����a���y�[���%���9����"	S�X���I�)�J��S��K�)��_��g����?u�9,�Qb�s�ǒ�%�*k�x�D��6�ٸ�����z���~2�����w� �9d.mS-�"���{b�Vu�����34a����&,ǂ)Ѐ���?�k57��?	�]1Xs<t�q�rϊݟ���/��x�6��h�;���Mm��(��>+;���r��KNN3C9�)��'�*�
lF�I�!�>����Q2qeUV��#V��+`�F�_���
���]��3w�(��|��������sNנ���l]��{d��i�BI�+w!E<:%=l��h+ROy ��\W�B�2��#��"�m��q����=#y0yEp,2ܽ�+�b�'~�.{&3�w�N�3��D���Ū����,ͣ�r�y�
'<�"����?�$�_b:�_s�q||?�C�+�yGg0�{r�.�_G��Ơk����~E���}��S^��L��i���ɾ_�\}U����p��n,�o�+^x/����ahJ�b3���F��"`������8�q�
���9��xi�PD'J��q�P$�<���FMC����"���S,��)s��Qr&���H�yx8'p�C�\"��g j\���<RH*�������!J/*���4�e���dk�ϙ;+R��H~5Ho��������:ʯ��f'�"cu$͊�w����L�G�n����#�y�5.:�>�@��:�ur94mo�W98#�'hx�M�v��v����N.,�'�7g���,�8�m$��=ợ��^ U�eO�H���z��h?��XG��2ㅘX�01���߻ocC(/�A^�X�\X��=#�?�w���(u�>{�Q̬?fٳ���A�?���>���Q7m�p)�x�!%��G
��B�SZ:������W���������4��Yg��ϫ6��ƛF׈^�p��
[ :��EG�J��\Ad�U8�~��m�ChA��-=�]�@��=zzҒ4C��̕t�M2��0����" ����_:g�,x���3�����9;�i�޳��Sˊ��;� ���q�P�q�g]b�������k��	�L�!vCp��Q���c Y�ghז�i�D8Io��V��ܴF�����j#�g̳>���q'����:9��A㟽�\f$`�>��I���NI���'l�pe<1Eh�^�[�o�x�.����침Z�!ĕbc�S湀�G�=���
臡�1����6Ww�{\�v��>���ʂ�=a�CI_W�ʽi}@�m�l�9��e�ު��W/��~Vu������t�(�.�5n�pj��[w.�}(8�u	�gɓ�r�������TZ�x�)>&H~pc��fV����`/�}Yw�k�w�r����u0�ޡ��\A0��f�.�]��/���6yS����-E�^{I�FƬoO���Ԡ��K=��hT,�~&�ץ��U߅,�+�a�m���a�z�+�eݩ��L<���s�+���j(�HZ�C�@H�Dޜ����oq������C���W�F��� �ާ��V�%][q�Y�"f��;�&F�Qy�ָn?,��� ���E6Й�6uK��)��?��-��aS����!G�D"s�����g;f!5�v�Q/�J���[���M�Y���ȻZ����J��&3R7}�B�	08�>�;m(�o0�I2�!}�{VB����|��LS�@_Űӯ�U��f#`�Ͼ���>�D��{�S��ȃ��}�,Š:�y�q�$��(����I����4���_�Ԋ�$�fӍG��_t])��*h���w�G'�z����� �)��A�R�#�g�	��naiل2t[ܪ�_Zq8�g+�_U���Ea�K�g{Tm����[g�W�;]������Yӯ���ͅ�������3T��R����T��K� BL?�$�V�K�G���FP/7�MFא�#���c��bU���?\�|��H��1_l�'��������lxg0�lӟ��l�2��+Kq,�D�X��w�u1���-Ǿ\�)���������X�5�]�AW~È��ݍ�R?]p��7�S��Zi���,UդD��NX����{"�\�t\pv-6�μ�>��n�����`6K���D��^i�9�F�y_����=j��k���_��m�������7Z/)̨�M>	�C��K��M�0A]m�<b�2|B4�!����ex]Mzn�>>c]���ah�5�0 �t��Gأ �Pa���P�3J =�%�����_-�׵Yy�W�A X+���!ho�T�Npʌ�㝰!�vL �o�+�ĥ�1P��f��� 9Y��ƹ��ȅC�O%�a|7�"�Z��Q��]D���桅��~E�tb;���|�9.k�̿�ч�ņ���~_D=��d}���a[M�L�0�z6����t���̭�������o	�p�sm����7���K��g�&MC�Kt��!+T��	jJc��T3%n~,��k�^��g!ؔ�s�T�;h�Q5w��ÿs���[sս�˾��/��Rz<��2���\�8{�nL�>��_d�U�y}t�GC�B!��k��̭�J�K�}��a�IoʦY�_��=� �������ͫ�2�U����V8
W�N���%p~>m��A���~��?#�^|7�+J�wJ��U��mBU���u.甄Q��h)3�v8ݽ����מ�UM
���}�N�䦔C�Ҝ0?�n	V�	��S�����~��Y�Тf�"�=c��S��V���a$�)��R�gc��|��w����C�k)Y�#γJW_S&�k%Y^�
)1���B��*� ����f
}��r�r���F֚�z�<,�d���oؗ�D�zV3���L��&���k��v���HBYiU�_w�(�aWt~����ҽ����ڋ	���+�FJ2�^	r3:K8f�4{BPջ��[9&���i3l%�Q���?��/���C�2;C<=�Ș�4pD�(��=�����tgW�#�����W-W�t[C�Ĭ���K�}G��F�[��>̢T��K��EĊ��2��AE����g�e�2Ӄ7^4~�_��F%�o��r�/(�q���hU��E�%ǭ� ��Gz�5��O����@�f�'���⥙"Lȯ�
b�qЂ���Sd#>�:d�B'�&�M^"h�=x�5�7�v��9C�D�L�å¦�Z��c��V��m(���|����Ao����^�|�\��(M���s�ǆ�,�����#\�{k��<�IQ��$��q��QQ��9F�}k�N@?�V������댢��Į��|IP��^��IO�u�&Iϐ����z�Vr��B� $�����W���M�^[$��vB�{1\g�?g��9�dp\��q
�3K�Dx%�%2������:4h�^����"9':"̄���k���M�Q�q�Oemv�"�&e�2p����l���We�5t�'(s��~��y�-��H�z��M��,�!'m���u��2ơ�n�R��J3���ԥ+��ʃv>�7+���n�;;LE�\*��ʮ�O����6�Rj~ї���ݗDf�܍�Q�&�4��^p�r�i�æW��'�w�7?>_*J�"O{�1�6��%�� 9AhF>W�QAv;O5�yQ}��ж\��/.gVʕ���"�������}��`$�\W�N[z�K�4Z�L���qHy�#�7A���{��ߎŬ�?Ԟ䉌o���NT�*��Yr��]C��$�ҏ�0NH�S=�#y�~>!��/���3(�Я2q�y0��p
ݶ��pw��^}�����Q0�s%�{	V>j��o���[E9o�Ы:��
��a��� /��4�������]Ik�s7�$����z����CG?Ƀ����v�V,�|X���5no7���D�a�im�ͪZ�����o|�wQ�!Y��dB��Y��~,'��#9���!���O9�#��㖽�$>�^��vП�x��h�8�$�VD���&j�y�������Ҟ[�|��٘Ģ:�Q�Ǖ��f�*������q�v�S��"��m%2�
M�b,%*�9�x�,_�� �G�����܄�xE%�3�Z=��N0��:�vCz��ts��jA0bm_�y.�u�Y]�\���7]����A�����CX��X�J����Џȉ4m��_Q��{iu�ye�;�'�~�v���{�K9�{?y��1?�/�t~S�:4�ƴ�d��q#A�����t�-
gsv/�Y���,�-{�DW��=M��YV ��:W�*䦻g����oP�q��M~��3t��-{�����طA����&����Ԭ�����?w{��]��s��Ikq��-,�o��\�Dw�Ԍ�E|��H���c��~�[�@�G�綢(�T?s�A@(�0�wgX����Aߖ�=��&u{y�2>N��{���ڮx�ǃ=�AV��lE���Zx��!_ӫ�}~�@�٥�N�W��	4�<7��5��d���4«�uo�0�-w�G`e}:��&��]�QM�C��y���㰙y��0�1ɑ�ɽ�ݩ��"�L'�?^�Hg���G����3`�&S���m�ؤ��L>��~U��_Z �n]	:\�i�s�|�HZ&'���[wQ�~^�޼Y��i��������ߎ��؆��VǾ��s<�a���w;I9tm�k�@�siRN��ۻ
�U<Y9����Bp���*���*�y���q��0��z{'��z�����E�T�����H(�Ƿ�u��}��~Z�F�`s�Nٳ/��U��=*�,�Ӓ�҄��~<��WL�G�.X"���l}W�>Ǩ%s�!�7��f���iP�k�?��x��������.[@i��z��6���H�]���<��,�x�y�����u��k��@l�E�&���q�oZ��c�uSW��X�+�Qg�`����\��3�L����j�vS<��7��>0�d��1�y�v>�,�<���v֘�^���;1q~\I����,5z��+t��K��
V�ۙL��XB�s��I�]�4��I}Y�r?���_������%�2�y��?Q�Od�=�v�K��)[�濵���I��g5�֐.X��4)�[(y㻭T(��=(}�%���Ÿ"㯏�ܩ;7�r/���)�V�2��	"�ju�}f`G^/�|��+c{�G:�,��`��G&�_�[QWǯ��}��;:�
s�{�J�S��3��s��Zm�J��mQ��%'�_VX�;���@��'��)��eF��ї<vy��tK��Q+9�xq�E��j#��]9ރ2\�J��뵛]8'�wL� ��F?ux95נue�Ǽ���e����f��/��lX���(g����@�f�J|�(K��q]ۤ���qe��3ZE�����ݰ��]����^\�Z4lW�8�赏�Uf��o���0e���j��E�ޠ��m@Ő�%�ǀ�Ti�:7���_�c��A��!�f�˩ιoSV�K#��{[��UMk�L���"������Ǚ�_����SP߾�Ln���Ȑ�7]���"�Y���s�������\y�f�f�g�]|�����������'�^�N򎷕���-|F)�i6��Zy�����'�^�q__q�T��(�����>�=� L(�^�O���j�(m˕gJ@+��
aӓ)�)q��^4���z�i5�L,����=���AA�$��b�u�#��e+�G�2h⢆���P�I��aW̺��a<�͙3����_E�q���7��Gy'2F%n����?�>��e>���r�N�6�	�E6���TC��
��ۡL����z�ۥ@�\	���?/�д%�-��8�3�o)Q�sB�:��KWFؤ�t�UL v~��H�A�?\�0�+��%W��>�;���Nh��[�`O�Q����..t��9x���]��
^|/Z�K�1�c;?��̙�5{�-�{f)<�V��Fw�t���f�O�e���WW~�\G�D杭���tT��|��v{��1v�3����2<��PØK�	V�!�z9�,�����t��7L:큾���g�K�� �� 4Ӷ�v�.���_r$�b�r���|>�)4�ݕ��;�Zv7���-=������F�vhUĻ��-�Q��>�f
3���TT�%g&��/��R�V�[Km2����%�v��&�l�a}_��n0�H��c�!�y��]M��.�`۴"%h�T��H���a��׵Kqo���A��Ӑe��7r�)������0׽�&�m������m��I��l+�����Փ�LSY�� �<�9�{�h�����y$n��z
�TOv��ݶ;�N�J׺�D�Q4:�U��x5�������P�%���o�vz���q���@����zl��!M�/g>��d��v�BAI�c*@s�����/��E�EBS��#eD�#c�K8����6�w�����*����i��?��������,��7Gԕ�O(%��~:���kx)KS��맼�:6��!�1 N%���ZS�#%P��EY��t��Ƕ0�aOP�kq�͹-r��\>�����5��]TRo̻-->f���~����x�}�U� �L�}�΅W�9� �i��7V:ٓ�Z�8;~�3�������N�@��fNTP���:���AȄ��fI��,�D�i/z�F
u�=b�N���TJ��)���޽���C+�C ��˵���~����3
��#�ߢ���}_f�v��w|A��m�E��7� ~6����o'��L��0i}K羪Îe3 jr(����+�|����N"�1
�F���N�����{~����Y������&F:��r��{�H�=�,&�l4�D�Ɓ!uE9;Lx6I��u��΅��w独?[ցe���
�nǶ��g>��%�;���c�����"**� ��#=��y���AT�sY���-ᕗ4+���z��J4!ԧ9!�u�j
���nwا��Z�U�����_l���'��إ9S�񷲔�R��sρ*e�s��b�k��wтb�k힖�q�kjr�9�4�}�E�E������(7�O��x�?��?Sd���P�4��Цx웴?&�{{�x��c��B(�a�	+<�Jc����.���g�k��
2����ڞ��9�nd]��~*�j�5:���vz-��~m��2�N
����\X���1��k����b���Zmy�ٴ��UX��R�k��iRݍc��JW��Hߡ�9�cK,���o�������r��倯�_�ViY�>Ú��Ѹ�3�;���I�"�/��[KYi�X��4��[��7�*�װ��vh�b}����`��A�2���u���y�����ՑY���;o���_{_5T%]��a��"����Ջ��|��
�	N�W߫	��� 'Xd}?W��r�4����s�� ov�d:�{�Yej�J5?3��cMp�Jݎ��t��B�$�N����b���J�Ӛ��?��2��tR�/kϪD:�����p�).���4՟k(taSһ��)R�ODe�-���9�������}��0M�D�d��؆��i�ah�ff�gGŧ��n���{W	ފ��~j�ެ1�x9��RM�>\���M�z(F'�}X«Xi��E�%P=�?&>SlYw� H�I�j[x��Ȝ�̕ꦱo�q��9���65��QCB*�����T���]2�����i����zG�
��>�
��0�C�]Q�#�r��v!��d(F�w��X�uE�ue�S�j�~	wn�:���FO��epJ�E��q(�b��� ~���#�](V�̟0u����`�?���m����Ԕ��`Q��A>�M��3	�E���Yr#�n-B5̸���)pe|x��h��Ҥ(H��ht�|�;C��Ea����4�P���P��PЭ�洵��K���6T�Q�j��-���J'M's�w%����n�hJ���џ:���j��eu1y��)h�2��M�U�E>��4��B�z|����{��vG����N=;Ct����@͇k?8�I����x/,q��i�9<���L�	/���~��*���TvE�T����U>��2�P��2j�aM�4>"���
w�YÞ��!�M�Z��"��|��[me|�&�[᣻=��/�M��ݣkh8z-.Ӎћ��?��}l�f�}Y��x�}2�B�Y|�T��Y�W�g1�"�89�t�2<;�+�u�^�`��9�1"LP�V�*�gO�����I����𷞎{E�R����v�ˡe�k������s�mY^n`~�V$����bC����ͬ��6��dM��H��������������r��-6z>M#��Qr��F�Qd������J�g�Ҧ��s�K��^�Ұ��J�<s�h�^R�o$�,���ө����4�k��a�*�����[�b��~���b�˟g��*�`X������� 󏒂Ф�^�w�z&���c�Q�LG��$��{Ĵ�S��z@'hf	�[{4,�	C96��3MO��vQ�Bs� l쬿F�0w�lH`�4D�4�㏉F��Q%�G��ٳ$<6�Eq��ХtPmL�����r�V�Pd��N�.�¤'eVhx]�:�oVBC
�l�2�y�+&�g{o��tv_�jsv0֊N�B���$Hl�t��jē��U.rZP-iv٣'2V8f-$�+�����FQ�f�9��jDA�f$����T�w�<�*�X��9��9E~��J\O���J!�����/�2u�Q������Ӳ���}jD)�������|+�+����Y j@B��	���YT�ݸ��6��tI���hB]��s�#N�V�&S+�~��*�!af����q=Hk\R�Յ3�������'�љ�� �/ݮ��;�ׇ�����AK1�f�R�	Ǒ�WO�E
��7OE1�v��&<�{�^����6�'GN+�0��t�^����[~+Eփ��K��~��:�����D[y���j�d~�Q88���i�=6����;i{*�����A����Pm�N����U���IJ�6��*��+S�g�#)ώR���{�(�(�.�@��eڴ�3��hJ4���l��V��du��%|��薱��Db� �������C���_BOm�?�x\�v��"ᶓq��όM������E��u�����cX������[��M�8��l9Oo��Hi���T��D�)��	&�
p�h}E]�j��F���/bld�]̵T���;��%Xú���N��6���`vû6D�Z�ⶵ#�&r�/��V�D���	�5cSg�n�*����+J�J�wQ����q6В��{�]�ö���5]��fl�/�]J���5��p��i3��m���~iMk��s+��C�ƪW���\�>{�i�V{t�U+H���<
p'c�	N�}��0[�;���H��~�"6& �
����0��<e�< Fbu5w)����[w���
����uB�ic@��,�|�!��5��uJo��t�J�fUD�ܮ[�b�Z��MCB�٧�e[͕w_?��l��p�f9��pr�70gi�:�[�<\䏦��s[�	 s�}$�������{������J��^(����~��Z�R���o*}�V:S�H�7}��-�Y����>>���A@���y �r���~)�r�{L�IG����L����K�+9;��AT��CkWw#��f���\�]	]�J�n�c\���}6�{aȩ�`����!��;b�T����@I	�3LW&�ϰ,��w4��٩1����������i�s��e���a����|S3(��Y"��*�n+�틭-���N&��J�ŝ���s�����Jۺ�:�YnK:Y��;+k2Yx#V}�'J*n[��t(���:��^lK�cK���S�9ٮ�f��(�}Sw�
t��k���M��Y8�㧠n�5�������g��[Y�!�뱜���b;e;d�#h�_]�9�mm��4��c�QS�� ��ݕ�����)�r	��6uu�!o5M��ޘ+țӷl�-��"�8?c�3s�:�M�H���ﻣI��c�e��A����~I�����_�Vg�`����]�3뮴���f�r�
%�0;���Ub�{cz�R��3�L���P�\� .n�	e^��& ���������o�ۆ�س�c�y�@1�UY�����������n���Ŵrs2����_���'�����Q#�p������f�[)(�sͩE�S^��&�����Ҡ���l$�B
��/����s!��V_W ���������bk�M��:���6
g�.�`��#���8����n,��x�&�{��/�
  �����#6�m"�*e�"9�m��O�|o�l��P�^�)�k���D�$R���)r�[�I,-��'�מ2xw����j�A^�}N-�Qa�=P�0�t	�d��������g0F��c��c�*�5M|*?����5w!Ř���w��x��{Q�q��K�Na���}����k���V����}�𰬛�zU؜^7Ve����O�ͼ���%�C�$���{}���#��&�;+^y2�xtb"ywW9�v��O��O��!{����	��~ڬ�/���/�����m���9�Ic����Х{���S�=�����Te��V��V�λ:��C[:�b%f#`�7��a%��Z	����ѹ�D<Y�(Y�
��M���; 9w�7C|#�{�-R������[ڴ��0�b;�偬ρ�
eN�h8	M�g��OGj}X���j��L^Ϭ��rK�g,s�p���w$7m��v	���J�_u��coD	5���O�d>��Q�S汹�>;&���I����}͝��*b9sɀ�}��~��$��F��^Z�Z�lE��X�64��)!�%5����+Qڏ����O����~w�L��=0��k��Y�yD܀�;5��-���
��cJ�j3(��o��ɐ���wk�Ȃ|!1��l_g�ϧ����}�T�rgF�4��lVS/qcg���+���X7�J�υ��g�օ>~�-%i�Ҳ�kϾ��~%B��!�	�B�����F�JrQ�'��7ɸ������tB������i)'��}���X�=�L����j��V���: �Q�I�5�q�{�'��������*���X�+k��ɬ��y�)�T�# :݌�� _���I ��Yͦ���>�&:Gw����_�k���6J :rm�����,+zo�S��.h���!�ԛ��
ƚo0�bg�^i�)�� 5�k�0�S���5\������b�������rcQּ����1=i� ��m�����n����-)?�q�4��F��'AuJ/�!�f�|R���o�X��7�m��^�J8��~��7z�_�Q�0i��?���[G%��j��z�Z�r=���z)�f�s������4��q1"$�,�5	o�VEN1dO�����@4}�e|��~�q�4���x�,.�>��J�K~[co�P��b%~1����� _^�u44�?�=ǹ���_��0zb��go�a����/|���Z?�{Y� f�^Ċנ(���s��Eύ�O���E�=EZ󩏗�J�Y��!�	Q)�']e�8�N�!w�^X��i��u��:V�S�F�G��3O�c��C�vJT�����Ll��۝�े�5���j>r���Hw;y�+��/��8�-\��E�CWYi7�#`^��(�8�%��}��{�a�n�q�X�7�����'���ؓ����dU?�ӓ=��y1�.�j~�^��%xu�Çz|{�D[x�P���k��x�nNڶ��[)����1��P�z1���6B_w��!��[N����T<V�ќ���X�G��Ɗؚ6y$�c@�����wm��ɦ�O_����=�.F��N�y�g!�{�L��<!�O�[��)~vn"{�x�{��������'���Z�O/��F���^�1ђbW��1�I��غ�x}��d���~]8�q�ܩ��;�aiz��ZY���urr���-A�-X]���Ig�Oz>�J�e�8�q͛"���d,�!CZ��1��Y����|�S��Ϋ
���YV��~�^�pJ.ӿ��%�����)8�Y�Sa�[<�"y@�c�QC��7b��	�qW;q��i5�س�W��� ���u*P^N`��s�Fs�6�>#\w-v�Tڂ3���z�:!�}���f&<4�s�G�c',<=��f�v�~���J���Z��$�]�����s�����l,�zH��b^\fP��Z�q8l��x"ۖu�ɯ�oU(W�bf�:H�T,��e&c�n�uJ�ɢ�x��
܉�w�K�<�\�D,���Mdٲ�r�� C���� ��s?7ݚ�X,����]�*����
�c��;��;M���!j�u�����)Ǟ������ڶAI�qGp�Or�<4�����e�Q�R��v�e]���WG�=�����琑�o2����mٓ/\��A4��D-��y��w�.�UuuXt��K�Y_��ɇ;I��u|���?Yu�z�X4�i��n�PN-�^iw���!�c���,R�2���،��a+�%���c��^���1e��Ѷ�eGN<}��br��Z����\��;E�{�ъ$ӕG���"�S��E�-������G,����17ç`�NS0wi�W�429g51Qw���϶7�zRf�� ����0��v�P/�ލP��h�"^z�Izd%`�r'i5K��~p(�����PN�9���ޅǓ�m�*����阬�t�%] գhݘX���:�������󫊄 �ؽ��س߿5����D�:�4��Ze*��]���8�c�}]G^���J��x�B�uJP<��/4e�¦S�@!� �Y������G:�
�ou��3hE2�}cj��)j��sd�ֶ;�2YB�Bh��;)�l�qv���{(���VD���q%��oV"hh�!���[P7B����@��UP^[�G>�eJ-��11�#�!PKM^:�?�d��tT�!#`���/�r����7r����e��p�ɾ�� k]��Lj�XN����c�8�d>P��4�Ε��܋{���bc�}�J�u%������{?~<Q�?��$�sq�rs��>6�n�V�~9vJ�y��/MD�Yt���*��nz��R\�*JZ���L��9O����x�ء Ld:����	z$y.,�	\x	K�RB�$\lY�ɪ֊`�:j�L9>b�6�&I��� � fe��U YuV���"7a��܁YJ-�X��6����['kdc��q��_��CW:��7�q>)݂�3,a��m"`A5'QGg ��U����E+�=�^CD��%� B�FF�FM� Q� �D1�(�{�2�����{&����χ�����{��^k����&���̝����D�wJ�*��G=��ƚ�)%y�L����h�&��MKV�I0�acƻ�Ԧ��~P4H�Px�Iww+�(QViM��u�O�[�ަ���;����&�<�ehz�Z���}|�@���J������c
>�b8�Vl�&̜ɚ�5/����a���à���f9�ώ���7E���?�k�*�xF���X|�:J�����ן�*�~ndFt�o�u�<H�}��nNn��U�w��5*F9�=z��z���50W��lJJ�4���C۝�M�m������^�� )�M�~�����\�ۦ1�UZu���N
s4$CgC9�3��M�虼�ɔL�#�o#$�{.�kBwCĠJ��^d�z�h/`x�y��5&�3Z�Ƴ�g��^:�\�y�Si��81�t�����t�h��.�,ވ�dy~��/W���@�Bq�F��E�6��/2>�͏�k����L��ZQ�4���@u���D^-�M�;�M�VՑ9x4S��7���
��t��ϽX��;jRQ���~k�S@~��8����SqIVzc[z��S�p���D���I�wΫ���R2z�e"�N��w���U����9�	U<�u�?�j�չ?� �X�9�3��%�	"U/���E_tQ��,R�U�^�'K��nI�k�����s��7Mk�ctn����`�8%������*0���%G]��;�U?&;+��&H���^�(��!b�{:���)�#�h�G���a�D�(kn�{����<>:����g��`q�4X��� �i�}@��k�
]_�PRK�u2�����s���&�e�u{�)�V�'}�mQa���C�*�(��:��f4`T&�A�7����!���)�s}�)u������p�䵶�';���0Z�a
��tV-S�K@�k�;�_�d���%4�"��[sv,+-k���ԭ��8��W�r��ь��H��v�aޚ^��#�-=�D��§�)&�ˌ�f�I��WQ�I��ɚ��h�~X�Ov����N7%�o��������??�������E�*�Y�ﯦ!�z�V��^���P��cY�@7M�(���j6���H�@|��u��2ì'��\
��Ƶ�o�02��f�$�T��ƶ����}_�[Q�x���~���N�᳓�O�;����i�PT��UZdZ�΀I�|���(ngH�z`� �>�
�M@�%`\�T�Ս�>
�W{��2B����^��7ފ�i�n�ɚ}�}Hm���}�=c�Hm6z�)�>��@���V�!j���)媊�Ŏ%�J��S�V�P� �сTm������i�s�ɭDթ2	�^����IHME����³�%�dH��gD���y+��V��*�&W��kϛ��yT��9�~X�4P����6{��fL�7��t�m�%6�95�@y[�^
�:L��/�C�����#s:�S�HN@�����B��yƪ52(��xh�t��7����Ҧ�|������>�`�{q�4�gX�"*L�|��@�6e��_�aѣ�T�T��'��x�7!��q6�ǡGv]i�XO���K}�c�V�{W�A�%z��[���o�JK��.@����ʱl ��R��=mz.���`}�k�*�nS�W!=f1����7�cv�5�)	r�V��/��<5�M�9R!�9�h���h����5po����8N��#�bZ�o`.�Ǘ���}襱6g���Pj�ց�>���	���;����<����N{{���T&~(ʫ�ѯ,2C�lpF���49�����Q,�X��Q֎	ǩ�4��^�K�=��
�W�h�*p�ϛz�����|i�M#�n�.F0����i��������X�<ӧ�~g,���O�)ƍ�m�iz����H?Gf���ɲR��j�ö�ߢ�?��ϙQ9r�n���:n�Z�;ëN�v�m��}x������_�F�ΰ��E9�䢤�~�l�ʺ]�?�|��ޜ:�c���7������1[�TH�0�7}4w�3ǆm���H���/v�,�V��v
�?��@�5��l>���\
?/��C�q��ö91F���52��3si�m��xS�Ў/0�����L|�V�x��p=�[��-����u_I�J!��\}�<��20��7o��L�;(*���t����r����m�5��9��Tn�)�<��;���17�������Ֆ�N�(�D�
�,�t�;�Y�^T���/Ɗ^�K_ELw�t7��>�����-����>����P��b�/�o����������r�:�A���bҽI�ߡ�}C��d(4�� ��!⽯��zZM�1��)q�����Y�o��v���+9T��D
{������,MJ��t���9�P�Z�,�bU�q�44U�$@0屇�Ԡʂ߇ r���R�r�{	ɍm �W���g]A��F��@8�l�zolE]�z+��C覎�LR��v1땹��FϻLP��;ݧӛ����P��
c%��YE�=J�zK�˛n�g��yZ����*����V�z��n�<ڈ8R��p?P�85V��uɦ��wBo������[O��_�X�4�`_��Kr�:��Ɵ�1����ӭ�ow��P~���in�+cX~���v��\&�͆, MwX�Z���Zy>/��e	$M�����:��N�; 3��)V��A�?N��WGM�b����q1{��#���`x7�Ńtf�a@�:O��mh���^Y}��"U��RV��iL.�_��5�S��������-.*Ldk ��;�b_������Y^ߋ�1N��
��ʳ�� �����e��/������<�bkkk��o�E���\��g�~�?�D�*���F9���s�.ƭ̺,pAO]N�,"�IىC��s0!��p�+��X�2�Z�Q˲h8�3�
�����WII��^���j��D��
�D��\4ZR_<�RR�H$J��p�g5]�)���Yh񼟭%]��%��8rw���:�Y�2����o�)j'��o���<6U��ͫ"��/v� =�~�V/�{�&������^�l5�~b�ؾiȟ���M=�w2�v-Z��*?��$��W�'om��e.H�N�]Ww�J�,ڣ���<�^���#�7E|�mME;����"������/��°o'VW����y��nJ^��̶]�i���X����\� ��e�'�K5��g�=V�5���J����������c	%��Q�e%_Ѐ��[W�P꫚�OR+��F�2�ţ2�j��l����T���K\��E'��)I��Z����T-h���gu[n^=�c�U�G��祺\�����PR�s��E�ξklxPl��鷽j
"�f�>����w5��B;4���"�z��w�v�a���Gd,�\�f*��B�'J[ge����S�^����^=SG�$����������Hw�D��r�
^����*�B�����qz�=�'us30! �ς������v�Jb�N`@�Q9k�9k_pn,�G���~U?�]]eG0(BڥT�a�S*�|?���TI[�X��#��a[��^U*�o�WW]V�������Kb��8c�N_V�B��j\H�Bb4R��c;-zӎ���8��U�Ŝ�,$���O���'oqw�1��z�NI��EM������2�S�F�Ѩ��R�Ţ�ڒ[���s�a�pK��� c�a}f�@@�u��$px�P��Q[�Q�9û����zeff� Ī��1��_���Ω(
d|x�3L���2��O��4I�:q���5���N��6��ym@wOV߽u�	g�1+�C4�:N2#���p�۔�G�aA�C#Vi�F%�����
e3;�9lX����|��`W1rJfPw<� �L�Mbw�3d�:�8w��C1�~ҿ��_cO�\�+��9b@�a�͞�҉��Yв�/��ؖ��td�O��^ת�e��L�0	�I�	�
F��{��C�H�nG����][m'GyݹI����^���ru��}j��_��ѩm�c��w��v�w�^yd�K�f�j�w�sO�Ы����������w>v�\"e�|��7��m�&�����7C+��Ss��~
���� ���������)��$�g���6��GY_p��xr�������퍅���0�b�N����~����3B�K�Sr�D��h+�Y+ �(H�>8�
6I��0E����q��!�!�w�5�σ
W���~��Oд_��?i_�z8<9���!�%�ɏ�s���S��6%A�;ga�zQ���'��NT�ԉ�S�Z�B�E``a����1�Eer�="���7S=8�C�.��ǣ'�t�|��`/֘w�2�3Zi�p�F��"����D�֯.�}Q�X��ۇ���d��f�8�K��򆷐î6��]]Crc�͋���,�pw��K�_S����$�H�J1�qx��С�ņ��I[B��A)�<���#��Ы�Qq�jN�>e���3���Zh�/Bo�֏O.�+V7R��+W���kX���?�:�$��,�u3����Xų����GeS+i�/s�Zc;M[���{��pS�R��"���kSb���eb��|��$:�4o�ݗ���TwTƧn�2ݧ� �3��|�勋�R�,Gv�ܳNJ��5^�Qu����O���˒���ǟ��纎�b���,��%�L��xށR֤��[�iq}���+�U�F�L��Ǟ�z}��١Q��9��x���@�7�ᖋ���R�&��O���+�`���o���{Í�}MlIk7�eo���W���3=�>l��j�R����$���ࠛ.�ݣQ���$=�H��͖qw��$��ҝ�{v��̅O��WYWON��'ҭ(5Ik�;� _�޻ݮ���^��&�N�J94���(�*�֧2����A���g���K�|΋h����R�a�L@ٳF���[꘸�~��!m���e� ��@���_,�@N�g�Y�@ϻJa�	\�<E?\^��Ն��Sٓ��y�H>�{���Kl�g�ύs>�j�h�>4����b��q#L�����!��g}}^=om��G�^�����J���x!��Rx/N�x3薛��?�~�u�q+Κ��&<�p���^2�K�4��`�\��q���;oh����xh��~_��nߏQ�N6x�F]>���d���0TCc!k$1#L���4,n˺��(��7z�i�>�8��_0�x3����o���?ʹ��IՕ*�O
^�5��C^��S�=��Z�g�����,HU��p�%Ds#S��r�i��4e'$J�σ��M=s" ��N���]�����/��n54���Ywj������-~jY�b�G*��k����8&,��7t�Ѱ���U�07m�DH��`ǫW���x����O�c~(�)�)$��#�E=�<�����dny����*��t���W=&�n,��;���m�K��J��]��P�c�FSj��x�Nfq���q�<�PLcԫ.��:T�{���y�阂�}G�f��.ˣ:�uxrb��:�SK��.*����1]�!���Gl�/-�Ɉ����Է���4_=}�x���k��ׇ�������>~ ~ֳ�K�J��pw��|PS�t�7|[%z�%tU���_���Cj��1�۵�Q��*������V��x�"�~�H�^z�T	&b�-�qe�����ۛ�O��︃i8}�>m':lh�Z���Ѫ\��#�7{���_#?6~�i�Y5�|w���?OA�ߍ�ٝ�� �����z�v�Cy#�������d����G�D�hm1*�_'iy���fn%�
����~����RG�����������b��d[pYG�'��"D��̚P��l��r�à5�j�@m
b='�Mњq:�x2�������6N�/Y�d�8�eQL�3m��_J�h�����u�9��1�An�/�"z׆]�ܨdS�b�����+�Y�/'�Z���~�2�3�OFX�%_lÆv�B5j)n��`Q���9��*��C��*����ƹۻ��o��_}�T��w�u����Y =�g1�7&z�k�Y��LԶ�P_�T�\g�cHAګ�����CL����I&. 4�+�-l�	�C����;;]�s[��m�/;\�{LyMV[L�1�х��Ҹ�H@���7*��f���Ύ�^G�-F̠�O�l=��y�CهV<C/�����_@�_��d�M����`�J�F,-`������v���fT,w�k:v�]�z�Yn]}#;�U�A��V���*�罡�R4��`�[]U'����1wLf�y�,�~Sj�d��r�D�	Uv�;�틑�����Ǝ�	���cW�<����!��r;O�v���������ͅ�t_�9�D� ���x:%M`��"�� �鹺13+�LW���VE�I=�R�����tw���M]mގ\��>�g���uI�Pؙo`���.b�� @�F���.(I�C~H9#�����;ث6��k�y��,ZInIu;��F��{w��#O{4��e3�"~�'�6���.;���V���6����C���oGgp����8�v&�y�<sv.��d����h���7��Z�^H�I��i�0�����|�Y��SS��֭��%��D��0go�(�h�mp"n�)C�;��gq��9޲����c`ǵ�3��
��I�Rn����3}��>��>@?TY����a�
�z�v�ŝ�'�� ܲ�r��_�	DY��6A��%ϟ��׹2�3v��qj�}�6����������Y8x
5��D�>0B
	`�����Z��"{��胁B��9�P��󉚜�ҁ�k���MnD��<8���:f���8
.c��^��:߾1�BɡC�H�J{4�=urN������W���4^���:C��3�Ѹ�1音|��,"Me~���ᢛf�?<;�1�LJB�����78��]/�b�\-9���Ͻ=w11/r��ҏBx/[{�_>{�S+ô�=5��VB��=f�g��z�,��ܙ!0P�&���I�
�t�dE�yh� H7��3�WPĄ:�z<�qХY>�'u�I�v1�/. 3���{��r����d�f�%f����n!�Ĵ���y-v���ot�tD%=(^���Q�ݳ����@*K����o�����\(�QjY�Q��V~�t6c3^'��#$Ww�F���7�Mﶴ�Ӭ9Ffgc�Β��$qXD nh�����4v��� �o�b�캊�ץ��L?�)	���Kÿ�|.�߻�h�m}:z�p·�S����}�4C\�q(����w�U�5dV�<�F9kؒ/��il��~Ӈ3J>��m� �E5g?
�K Cw��5d�X%�������2	�����0E��|[-c��Z`�?���1�8�2����u�W�{j/2�[.���ʁIUė�F^�����*�!H�(J���ˮR�>��f���0KO�Ң��D��-��6��=�fKR�0�w�&ˬ�����;M���^sn���Nk���h#F6�o�w��k�rU�鶘F����e5{��Yѿ!�5����>L�Ԍ뵆�s��<J�@)��)���Fe8_�}������������~�f���O�d'�,������Ɲ ����˘�b�˝G?�)�y��_��t�J�nT�s����W�
5��J�7G�:��p\X%ޯʗ�|��v�ˌ\/��="#L@A��������I'B�[j�)�0�x���Mu��(�}fh�dH�����ճ�)���ȝc��b��嗗�2�@r�~�a� nM���8��0w���n����r��9�)GG3�0}��ɏ��.|Q��`Wa�Jm�( ���	7V���h�r���K?�0��侜2���j�HΝ�7��Ư`�h�j��P�0��9AZB���rR�K�䐷*�US�~���|O��/��pU���FT4�9Ŧ�P�BL���5�l�{����ҳ�p]�	��n�ʒ_��N(%j������l�;�?�_>���&��ͽ�nx8.{t���.A��q��m�HdրZ���,9{�yrʐ�"�ɨ��	�L�l�a��-SF	����p��!�㊪o$����7���a�E��NR��,��B~�����;D�> o;N�(�۔� ��k����]�n/�
CkX�.$�]x��U{�Q�_O�y��9���h��0X,�Z5Z������;��U�?����yG�*�,����d���gF�@�VVB���f�ym�g2|�<X"���[�#���D��R�]������&�z�O�z�:��`��Pw�׏�z�?�$�, �����kۓ�ma���0�3��k%�bF�E�(�er�gv[�$u�ۦAy]߫avO	a��m�]ZK�ky����7U�R�1�h�K�UTV��������k�#�C�Gq����5�� lA~��ks@)nsՕb3�p���8����������p�����5��Iw?��0٥#��@洅D�Z��c�����ӈ0�V9���΁�@�ߺZ�\D�=�������1P��MIz��{��'��9�x�tҩa?��ۥa��S�ž+�rʣ����H��S�Tr�f���qP^�3ɏ~qţr��C�\�l��(�3* Ҳ@�Q���t�LXj�;H譟��cc�q`�s��x3�U�m6_o����J>k���RD�Ĭ�|�[m�w�-b2���I�o�-�hg���>�yկ'�TB��%��W�lw[O1{,~��y��\!���� hbݪ�WPJL� ��K�ڀ3Vپ���R�/��6�M���p��<ڀ�g��<�C�����ն�Cnv�%��k& O�khqXY��� <�'{��˓�i��8٧즌2��߼�^�(Ơ����"�o�&���l������Z�\X�BCƸ��3��&VP�-�!���WoU���.3ɅXN�y�M%*ՠ�o<"Aޟ����,]!ȧMQOS5��ȳA5��8q����UUc �����;���e��j���d�	��7�")�Sb��?����֑Z�s?�=P�N�#�2��)5>�������aI���F�Ib�s��t�*Jr��n�!�P���^<���M
N�=����۟�6�4�RBL��Ef�y�Z�x/�o��L��3F*�:5_y�Y�t��A�.�	*�Z�Jo��\Γ�67�'�H;�u�w$@�M)���JP�D�������<Mat�?�_��0^#,�É0mGOC>�n�3�n�W�3��o� T��[Gmjſ�sUʇ�xks7�8/Ԧ�U�����I����������<'%���_�I届ij���}�t(��Փ�)}��e��f}jy33&��l�3����Gܐ _i~���b4Rt��F���Gc샼�[BR�v1���-�O��QcѨ�-��6�u�%x^��w��տʣM�U�����o%���N��;�����Q�ڹA	nzm31I˥�o���fJ�<��y�K{��#uu>�ɦ%_�_���N9wl#a I�Ҥ��H���d�5T0��@쉕��^߬���5����i���6�D��lu��I��hS��A��)� ,;^�~�{3�ЎO|P�ǆ���( 7t�N��� ����T�x�q���Gf���x�(_���%�J@���b�U3���� ���G��9L]!���E��Uo��-����s��J��_�Ï2��+�p/��;Y"���٦�j0%'���`s��xw)���,Q)��֛P��Z/�豯�̢���e�z�@Z/X�bߦb�]6E�t�c�M�j$�=��Xiܓ<�R�M�{�ak7�x����5���d�-����zO���(x��X�o��1�l��O�R`&ݕ|�*�z��+ȝ�]^��*@����{�̧�����e��5��~�H�q#I��a����*�\Ed�SP��f�p#�5*MH���J�h��4u�C*V��|�&�N���$��dd||��ӟx�������g��2;;`���V$jOn6��_�ƾ-X ��11S���[!-9G�\?�#�y����i�Ɣ�wP]!����'zo�]�����An�>d�ߍrT�~%�����`L�c��Ph7���06�I_P��f:h(���M����eP�΋�
895E���"�G�8E��H%�T��'��;>]�.� gv��l]喞�����>y�v�D����vV�#O�'XUՌ���^5a�h��1Q>o�3웯^��q] ��= o�˓�(��7�)(Fnhǂ5L�-��>��:\[������	������"��`GX��F�����C��VM���]�
VV9L�I?�M�u�b����i�����=I�1�ПJ2�d�͚gw�Ԟ��F.�-�x�qK�N��nE�O�К�.��~�o��vɋ<+��_R��rU�����E(tL�l앾~T�����C*�*d 8��Ch������O��]�Xf3��5��W2XO�����_F���.�nTC�|n^==`Ԩe&�#ii�wh���Bܬ�v��Yu߭���O��sN4�����h)�Â ��=�%{��!�O�x]��B�� ��mn����U�wH�!�5��ܔ��$�X�x���Q�fV�5�V0��W��
v0K�=�6?�ٜ-�q�(B��l�B����,�R���7:��v����T�H%Q(��R��0�	�|hk����tk��j�:�d�5M�b�~e9�,���8�8��]�%���4b�ޚ��3xA�;1�t��E�^����e�_ =VgRz6���� �Дi��I�r�w'�8�w���D�d��Rɀӗ��J}�Jp�8���J�=]�X���q]c�x%��uW`T�G�Jv�� �i���q���*fXkƵ������Ų0M}���uc���ٮ��t���*�Y��
/��5�z�������}.�m������)N����/�|:���I�aO��:"ט߮��|Yv\���W�Gw�z5��w�S���+Ot ��d��[u��\��@;Y��tx��Ʒ�sSl�\W�;�����|͖�2G|���B��PR�oo���zlll�9�yN3-j�9Kь'"dh�mh�3���HR��D��<֩�s7��6�#�S��͏��cM'��v?��S���^�AE%W>A,��
a�<�R���6�^��*Ӽ�eO��Y!w��L�x�׫�;ְ;wLк����{��t��8�&;����(�.c���|[`�w(ĽP����EE�HH.
���ny
���xQ'Hc���kf#[xoN���S�1�󱃈���C2ҭO���&�D����6W��3�u�|����_ً��D��m\4�Y�&_��FΜ�u��nb�~��e���DO��W��_�G��k�IzF�7�{I����JM����Z>��F{��C�U�5^�����?*.���hݡ�URR�eo	�-G�*, ;k3��Q��(���j�Q��S�ta�z����D@�m�����"=�b�ѓ�f��S%���\1��1�,�q�.�-����jH|���ꪄ� �j^�W�g[�u�x�Y48��
���[�l5Vj�����ފ}��-M���]�L1ٰ�擡O(��m�w|G�Ff_r�'���o{Y��6b�00Iʫ�NNF] ��#�G1�/ƂU=�,<��$�1
�:{F�n��fyQ����WDd�,��i��}6U��D��΢'Y�X�d�K�|��19V�֕o��VDщ�:=��%
e��9�8_knZ5k6&h*.&nI��H]y�8'���7 ���O����h��ŋ���O�}#|�6�A����ǀnY~t�E�/I{�K t�i@)��L8&������M�߶@���ޛ�9C�Y���x��#W�7�)��\�i�qj���-	��o��Y�7Mֶ6�q��ƲD������0ܡ��cO7�*��1	V˥�w�K��j��Z��0�ޔe,Z ���� {�^��6�FJ��I��ɜYl�
7����ok��)����p��>]��{��syTΓG�k8�^q����Yi���:7�d~��:�����ڟ��R�HI�o�wW�uo)���j+�r���*
� ���EJ�Z�4�+����>��y͖�y��mSB��{���>#
E-�[��8JH�x�U{���m �Can.v���	���)y�n5�);�����zY��Q�	�k+�[p����Ǔ���D@
�����Nem)5ad�LY��	7�*�.%�xa������e�ݠ��E��Ek�[�D���ԻSRN�pS����Ɍ,�qv�)h� �,O9W
��!�s��n����U��/m���m��	Y&m���Ť\0�?�z�'��"!N;8R�Y���s�!?X�[`39070L&]�G9�-H!j�=�n�S$~�n�^���Gg;m�WO�A�}P���z��d�W\p�/��m�Lc��umꌗ��<�!��fX�`�����
OM��(�Ռ��L���V�!�l��+����/�A�0�n�jzu�#�'�"3��<U�OB��U���*:D��ϛ2�c``@#��}U�9�=p����Q��:%=`clN�w�0Hn<�~ qBJ��"��kՎG%w����K�mE`a"��͐�㆛3�E�Ѥ�:���l����R��+{�3�I1��.���)ӑ<��P���Q7g�7_�x�q��[�re\*����c_7��
(���M���q_�B8ߐ�D�a�tĤ���v��f�E��n�KѤ8�m/����+��y�d�$��=��)�@��w~��b�l<�5ZW��v�\8�,�jy�� I�9w���7y�k�j�O-W<x}��;|�!��e%>Ɠ���:ш�,SWl��ݞ��S�ǚ��:5zx��_�

w�|���JWo`Y��p�5�E+@it�k��q#2���9X�U���S���+[�oZ�~� ��Ksp�3C#�-��-�N��]wf��X����R&b�M}0�5ވ�T���w.�\M�����8;�O>P��0Y�1�!�z��xi�B��U��[�{�QO�K�_F7��$L����%��2+��
����T�η���K���<��heԆw���΅����7��/�o�	Ҳu�Lh���ͭDW`O�#��%&P��Re��! ��%pp^0Ĉ3/A��]��p��M�{�!U7���O��1%���BggM��O��JDm?)^JUΨG�"�(�g�J\D���:��#ݦ'������>mt.��yZ��9R�uU�49|���lN�2�!T�������va,y93�r��;<���#�e�� ]�� �����S��lE*�:g
M�u�W�Vvz�jA˽:��(�r�Pm��a��jh"(%C3�m� ��v�ҝM��y���H���z�Ѹ�0����)�+��,Y冊�+?�yB��:z&�+L�؏�a��-+��!�������̑���ᱱw�;�C��<T��H:���۳o�Meu�*�OD=h^?ư��6���~�N4��?>���g���{�E���
�Zϔ�^-Y�|Asa;��K<��,M��8�z_W��Q�Ե]*Y�e2�o�R!��w�#6��ւ9�:�U'&��ŷ��Jؠ�4ژ߿��N}&,L�5����Z�H�y��FI�Bꣾ Co����[�i?.���$�����H�N][[�g�7S����%��
!��`���:�6��N� -�Ȋf�ObZ��8�kG�9VD=?�Wt{�+���9�q}-D�ҒZU��^ɔ_�
��b��U��f�o��ԛ���Hg�YV����ɾ�t���Q�zrOqYb	����^�96��7 �Ặ����K�eLMt�����K�9I^ܗ�W­���~0��Ճ��d#��1R|GG�ڋmXv17�iÚ���v�7�o�%E��������(�%�|V�-$���D�0����wEM3�����O�wtV��i�^�qGY�ɫ�:����:���T��5"Tf��ZVC��R�?r,I��3�qo�y5���۶�^ ޒ�%~I͡q�i�9�ף�ພu2�K/3"�c,�l����m{A�GQgL�R��# nBS�i|�=O��D"������rx!����s]e
r�F�a\
�Zۇ�뚶�H�*�3�y}K��Bf�R�(��s�-�X��Q��J����7f��n���'"���{
�K�ȫe[��`�`�z����P��C�Y�y�f��z_�u�c	��j:C�b-�|4�8V����'U"Zc��7�����0+�6Z�W;��;&;~Ԕ�{��Q���lb.���
\N��`�Ɋ�J�d���"���/z�|sŪ3�SS�yj�L�=�:n��b�����L��IG!0�������a��,Y�q�G���Ø!����g�����_Z��n#M�J��H����K&����z�'M�B��I+����1�����j��2q�妙#<���xݫ��ZW�W�;�&3�v�IE���I`cc�\�uU:L�5�~�86�{�j����`��;�3������a�&~���[��IY��Ϲ��?�T��}���]_f�j����IU<僜Z�*��B��'f���نG�V޻몵6.-o��' *)��j�f�8�Q�������e��aj'^���U��A)� Ą���"X*��{�+��Y�L��@��ܲo�b����	��a�A�^B��/v�:�\tϺ�/�] @u�L�z���6 �]��wZI�55�����a��:\y<�ZL�ۮ4��T�嘐|��Q#��͢�RO���c��gxnܨ����ژKGT��̶��vu,��G�>M<���G>�kó�D^�oH˱v�I%վ��-�o���V�k�q���HA3ǫi�؊��%��O����f3�U-��^g~�l�+3���0�П�+j��\&Eo�9W]v�XƎ���K	�H������H�^�=Ɛ�ۚ���g��Xa���U̯Oy1/��}�D5}����#����B�u]�u��m%�Zx�u��Ο�F鼗�>u��:�s��tx����p�����[�J�!��!�c=<Q�z`���a�.^\W��C����y�a��g'ޯf0PA��D�����v���rd�"�㌮J�k�gY݁(¼�f�X�}<F�ߘ�����L0q�Fw�ثZph+R���a���t�@�(��{܉r�X$̛����޾�F'��_�7�N�ԫ�����0�b�	�Q�����m�cK�Ep�����m|F N����z�������Z[�^�� �ICl��	�^�OC�8�M@��93����ZYWJ�\�M�9�O$�ʗ�OC���\�7�?7��`0�&� 
��,u�l���TE�,M��9��j����f��P�����# 9=6U��5�(=�{���G?0fD n�"?��e��|���p�_�����E�'L�eGY-�v���*z�yE�����.,1Y^ԣ�Ƃ&2<�o	���!^͖dh{�Y4+�L����ђ>��`j��_{����#�~]G�E�ryҜ���,�!|E^'�J�A�}�b%Wl���]�Yϊ��{�ġ|��lQ�\��.Mu5MA� ��?qe���K��mm�ޕ�lwĳ)]~x�W�򔸐D���F���1.dgDF�3�����u�s��
��4�(��~nH�<��{ү7����H�!��'F\w� m��yo0g���|zl�[hT�fO��y�7#s_Sy�D�i�Ϛ��Y�dC�Y��d"J<�+Z	4>��ȇU7A%T(u�8U`�xF�gJ��t��T9r��q.�)�#�@߮{ygҴO1�.u����J�s�b�,���*�^��m�x�L���^�_Q`���ғ>������n��*�P�_d� MB���5��尃$��-�m�\��^��˚1��G$RY"*����m��cR�r5����>�F�����������ms��(��|���YS9��{��BRQ#ToX��w���3ȶu[����T����hrF��C�����yf`���Ԝ�y�ӭ�&?0x/�$ ��,���&�������CI�Գ���FN"s�<==�|�#����~&�抋����v_R},�!U�bob&���䑼\�h@�F��v�xw�������$9�U5�v��-C+�Ku�h_Pu�ؾ��k��^يqBF�Q��tK�P�/��һ��'���|Ax49�ƛ�P;6�/c0M^i\�4��i5/ݢ携V���>����6S~+�9��/����t�2�\PGĊ7��<����F�oh����O��d��VҖ�x��cb�g��H<�p8ܠ���]{�h8S��w�.ҧ����Y����ޣ��wܲ� Ld��4޵3��)��0�O	�h������5&F.Q�Kx���.�Ў��/4nO�ԑ�[���n���v#�y��U�Gh&�Y��[�eN�1㚿������p���V�u
�lzr>;z��^��N�4%5N�����]v�B�	(��%�;<0�`�P\&Ҩ��"��DDD����%��¡�2;�y-��'峺_��<�#�W��w,�����nH20L��.@��D�Ueq�#�,\���dA��������/�?_�u�R$}|�أ��j0ʈ;�E/����j�T�c$48����E�:�ڣ��	�3�\�&���\�
[%9�Ӕ�[r����}��	ͫ8$�����t>��V�")������3�.'D���'ۆ��R����{�e #�w5F�ȏ��,߸E��=_���IQ�X�)i*����3m�I��u�Ѩ��7"!�kbu�X�5��}I*t�Ru�gy��غn��99�&���P����"Z�X�I�,ϻ�,q;bN-�/��zn����e�q?^+��[�o���^�lmA�&Q�7�w�\w�n���Y�X�C�@�� @@�?���ͮi���݊�S\JCqi���S ���V�ŵhq�ܵ8	V��]��y�极�C����ڹK~��3'�.�ee���U�B|����*���������1o7KAU�+��Q�SJ��0�g�.�?X����[	�x	^^���q�^�=�z"�
)s�q^�� j~KU��d��Y(�9/��:ܭTX��0�R�E����{�Uj|�Z�LTr�m����Nʹ�ҧ[6n�Tg6�'I�s��_BL���>`�O�o���")n�J��MMH;,}�`�̋Wk1E��EMN�,�e�J�YV���7;AB�x�V��~��==�_Nru��@#�p 1��O�f:��'}�l��TP�
�[��������$Y�I�ϒ�x�ە��A��D�"���ӗ�$UaE�����}v��O�}g«7���H��_�T��GƶZ��^ �ˤN6~��������@��ab�'q~5��D}�.�A�ĳ⮡�XB�w��@����X>�ήK����!���T������g9p:j�;K���Ӑ����g��������wpd�!�ǌ�	8}\�����_m~��(�H���[	&�;*�~ES���ߜ�ߐ�+�t��,Ѵ1o��ꑀ�d[��z��qWsۦ�6�ZYjeȋĪ�zaT�Nw"��W^{Q�Uۛx�dk�U{�<Fh�����PM��N�`��hU�d�_\Gk��(`�gy��A�R��0v6�կ����Ը�h�{tt)AX�%��ws�4�RB��QHK��JR��Y��o"�!F&5drR�v���i��+5�l��C;��/�=MA�D���q�׬"��U���=+r�P��r���2���O��p�j�W(a��3iz��	ڛ'�i^x�8n������D%J�.���)�rR��Xկ����|^���4�O��
��R��M�Дy��K}�N/A롨�ٙ�y��ll�~u��=���J)nx��A�e��?+�XA�#���v�ŮX1��y�z�������ګ����T��cQ��(u���d#	\�ՆT}�j����l�3�b���P���6��ͫOj`�F'�CP���>=��dX.��o��f,̩��&�䴵���o�W�3�_�%���B��	�s�|K/ ���g�M�y�����	�O;i�g�o��j2�c�]5@�<X׮:�66"_^!��h
j��oA�]�z=b<�92 ��nұ��z*���@,�3�#��E#�(N3�]�')�',��w�_%0�Z�>-�뭇��?T����Al�����y�Wf��4PE��G��,yt��,��H����{�ɅL����6b����udKXH�tߧ�X�=/��LOU�w �Mz���[����7��""ˁ{7��A˿b�}�^��C+��>��~���pd��8�ɫ�#����r��Gx����ڰ���a�ƴ�%.����k�%�-՚]w&<�����Iu5i�r��K���j����-�\�n{B���fӢI�F_$�<�NF��aSv7��d���N3cBK �;O�13�_mv��du���i���Pu���R��Gn�ƪ6�ƮnR#��52t5���f\b�q��9/1�o������#_��Px��s�1��������2�sv�9�2�<9MN)�z�{�M#��A�c#��]����ě�?8�V{��F�V���*_�nB������q(��]���g�6�8I�s[�Х���� �`�V��A��N۸\v2\��qZi%(/g ��Yԯz��#g����r����F����lD���[�Й�Jr-c����FC�(�OD��ԅ �2���Q����#7c>]��mo�.>C���l_vP���Se�ǭ#�O�݅�^?`���z����NQw�\�� ��:���O��Q1UG��@�te�U!Ѕ�B'oG�=O��=�9�����7;S�D;�];����������a�Pd�!K�9���m�N/"�[��ZH�'�-�S�^[�x��9������5�����b����������.+Q�7_�6^jv�
���=�-�We��ۄ�e��BM��O�2����_�`��a�*"�;^�y	�Η�f�&ݖؘ}���}V~/���g^�V���e��+�a���:�����L9�(��g.�|��#�g^,b�E�
B�'3/+ս��p�����g�����DG�5"�F��K��!�	[dՓDS�ry��x`4�J�ޫ�ax� �'mS��p�~V�>>��h"V��{_�d�POe��� ��F�HZ�{}������+����� ���s@݀j�g���U1J%��;���{;�����e�J������c�|�	f���"���9o���%�X.WqԃI}�ڇd��o�i�����b�������L���u�$T���~��q6N���JF#��7#�o�}�ȪAG�uԐPݾ��Řd]���O��#��F��<�A�h�?!�jN^��ۋ��g*o��l��熃ߩ`>Gk݌�u^F����ۃ:�����G߶����8�A���q��{�d�H܁���4����, n��U�*5V�"J�M~k�Z38\���AB���H�3�)k��3R���pe���c�2c��~y^��YVň8&�Lˍ5����H���Y	��=��ŵ�؃�V�H[\���k�����f����u��������||!��{*�{{'X�2e��

8/�i���'�D�3 r3�p�tԟ�KԲR�
Ӵ�Q��$C�&!m���Џ�<�^1����~�~�xL�pQ{�M��
�<G��w����[�ʇ��C	!y�H�Y7��wC���S=?�
)m�1�����u*�~F���b�L��A��nF���d,�M:ƭ����ȞL>jk��}�x�,,,�N|�=xS��y��j{�i��+��虑4}�7�Y�as�����+��?_�i����z�̼g"����*�/jhK�XC��;�)��N�B �^��N�A�ښ	"�vu�F�!X�G\,nՏ��������S<{���>��D��1 �c�U!��-DG���[9МJ+(�sk����s�LKG<r
�p<�����Zg)6�j�-Nt~~���
�6�D�J��h�����`*��d�Yxt�}��II��j��6HS���OĉВX'�z 5"@���IBJ*�M4N�+�=�����r�	lzex��:���r4���ٔ.׮�?W�<i	�k�m\�/�q�4`
`ꬷ����x�ڍ 	�̰�N�󋋍L�jwjK�8�7�Z���䊥�%�_d��U	�B)m���~Y.6�(�{�.�f���3?����?�$l�hjl�R@���B�V�R*�����Ŀ�y��iV���)�/L����ȳ���i${C�䄳��7�P�YgV�l�=��;K(x�>l��mӦ%̽�]��}O��$a"לF[WD��M]��)�ݵ�8�����iG���n7��k�gY�9myy�4I��O�L{�o����9:�"r�v�f�~M&薕^�����
�@A����&����71�2 3�I5��sZ�{ā�9kS��O���xm�K���j�T�u���9�0�F���Dp̄��<mH���C�9`mwiCؕ�6��{fc��k�%�B�\Xc�O��% 
]����魆l��)
�T/K�Zv7���1E�>E���6��9Η��y����ڔ��T����u�ZM��P:�������z�8�^tJ�Ȏz�(2Xj�����Q�0�BP�� �d���ܸ舋�C�����[���efy�1��0�/�8��aO\��V���ʐL�&ǜ'�.)5��n��h�bS�);�ro\������ۘm�� �A��E}pҕ�R�ep�v7~+s+n��E�����Ĕᖮg\�[�>ΩgKp�(�nk��4?L	�aw���RɎ����~�A����[v��o������)��qωe#K>��T#��
u��u$˫��޳IG�&T��_u�����y�A�~ü�k֐�ĸ���Ĕ�s�tZHk����2�����f;���Aۭ�b��\��eX<	l�X��6�e�����S�Hl��W����Z�G��m}6 �X�5���x�h��m�DT��� �>��9����.*N�;V'���b#�p%+kT� %��I�Ml�[gD�&ݜA._���:��O�{~�˥L��<��f���t�~�e�%�6�Jq����zҘ�lW����m��U�Ɨ����jS���S���ҋdۺ�\��)Sᨂ�6L�|
��'�N���}�r�sX���,���E;p�|��F��P�B���[���B �^��M�I`�ː�e%W�i���ճ5�Gx8�A�0�	z�S��L륚�	G���e�zxԓi�~�CV���E#6���ۗ�N&�6�Z.s��s���p�|u�_p"�$nUV��r�w*��Wow��m�%�Y����˴!�k*;	��O�Lټ��5i[�dj���*<��fKQ¾:�ZC\��� %����C�i�| ���"������Y
���t���(2��?.��k 	`���ƿ^��Z+�����R�fk�?��no��ı���]G�F0�D�A�ƴ�~�}|����|���٩�ZY���cԊ�JU1�'�[��13d�U�vY��^��>@K�\L�m�c��h��K�<��I/�3~��4B��'�Z�<��1�;�7;����n��cuC����L�cy;w��]�γuM�~�Dv��Dni�#���W+�o��.�m���oO-˗Q۷"czs���گ�311r���Ai_�c����I�j^c�D����`aqg�0Q)茍�`�ض�(�l�}��Ôp`<�aHP;]Rg�]��lx�����#�k�J�5�4�"2NHU�?�Ѫ�U_��b^Ub�*���S?�N?��v�r��G!�͍LL������D۾����^%t�"�� �'R5R�S�Bf�;��^�s�}>Y�����41����6"����-�dU:�ǝ���@<�'���6M�OY�_k�e�(��
��ǰ�T���@���C> JD9�}�����N���z��gJ�%W�r�~�&A��:�xd���!�i��'���V'F�f��S�/x�O+u���*/�?7��|�T�-�d#���H'��v�ګ��R{�Tm�l�@ʫ<(��8<��9���=�ݞ��8q(�T����M9e�����!W�7��8i�#fǃ�6�{~a�Y��"6�K�ΕW}2y��9B�al�Pp�nΧW�R�4����[�����f��Nl�}�~�eOm-_���6�t�(�R�~��}I!��;vNU���߂\���őD�{�@���uM��i��-e�߳�����1Ѝ���ظ�;S���GJ����Q��K�r����9�ҝ�e.$ѓ�U)qp��4�vN%<��,)�"������h�L%��uz7y�m��`�`�_C�f^b���Fm'�PG�gD�B���9�)��ׂB߻F����P`\N�ާŵ�d��}&�D�/c��פ�dk.O=�8��Q/�|V�WJ=%a���UJ��o���������\�k���B �Ͽ�Z=��"��i��0	Uuu�$E3䆜}���,�S�E��n�\9*Ȯ�ҩ&�$�ʎ0Ɯ�SW�,D�lv/<�����Z0譊���z��LH�q0S͌�?���������f����z����bv����L)1��h˫l�	�V�����\).��3��r�q�W�6ږ)h�?�ʿ���i�l^��T�v���w�m=}�}�i��Bhi��X`l�M(w�Ӎ*y1�4��Ŷ"@���#>Iɸ�#�:�������6_S��c)z��f��/���<��ue���&.bEYY kX�_+3ee�v���P��s��� �{�I�m.)^���f"ޜ�א@e���� r�6���b�ۣ��W�"�c*�k�|D���U�۵�TB��t��+���i����,^��f(�ߥV��6�\>��
��d�?�	[XV.�O`�[GDF�\�� �����71�����{o�٧Fجb����̷�/#�8aevi>r��vN�=��k�B����7DCz�?���pc>�����W��
K?L�����t����O�ǲ�'���/���\�-�0�)���-:X�;ݹT�t�~��,�f�q$�m��B�D���/�R/�������[����%���V��L�i0l�#�@�㰕@��� h�_�������va����YEs��ʁA+�K'�>+[BT��rΏ�/2�eH����2x0xڵ���I���S+�Ab�eDp���1�]š7&�'Ϥ��}��(�Iʱ������fܮ- �Iw�)����'ө=�){=�nD����x���ɼ|ʷᚍv-j����Ck�hu��@�i����F��ْK�O��a�[��['��Z��r�������#~)޹OߛtW��J�+h0�1��Fޠ}�¥��z���K���sK$�*�Xtc5{�o��qew���g�}�HJ�
����(�.ϯ^��,�L��x�5t����,<<��J|gmPN�
8��w����.�@#s*�%b����B?�~�30��Ya[����Ѡ$3�l�E�/;��O�J��F&�Y6F��k9�-НR_X�+6@�b���;y�Yμu)[ŌVP~(��ݣ@I��<�HA�I��'*>n��iH��-Iv�g�!����1=�S����O҃vS]����hy[����DR�R��ˑ�6��c5�ӯ�1�|�H�yFi��F�^�p'	�'��Q�j�.;4��bn9����n2����� E���׍�Q�2��g">:�#H�KKli����/+�hE���B��s\����1	7���Me	���1vx�^��?���X�0}�2�TJO����B�[�f�Q�6_��ч�Ē���Vnn�2Sw`���n�b	'wl\��U6j����6�C���K�tC1b��"�?���f\2���r�9��dL��%�+�l�FQr'��q�OQ�~й��s�z~g�m�v����)Ns���?����<R �m�qCbʧ9�}��#R@W�٬��VQ��*6�[a�<\,��M�V�R���vX�\{V���ɍ��@X"aƟ�A备 �Iaq�t'5��b[���@��P�-���ܠ����7q����	�o9�}^�O+\0=
H���s��qs��|�s�ы�6p]�I����'����V��G�VR[�v�OI�����|52X�b��o���]�U��̄)}�1�'�6���5�W���2�vÛ�a�07�T���ƶD�^��ߋT��yF�5�(�T��m�����͈�v�)���HխA�o�U|`3J�`O4G�˻�~���.%"���]��7��^������X=��;в���oq�f�3��2��}p���(~��	��*�Rּ숈Ӣ.
?P��ԫ�Xf�*�U·�W��Ry$���昕�L�_ ��Bg���t�f���bײ|}�����E�(��aqܳ��+��@�?7�e�dRe�j�zٴ#vJ͎��)30�$X��!?�'��u=cod_C�D8��f8�����O��wlmm�q���lj�e'��K ��v���=�2��b��Y�=�a�p�BG?��0�|�lw��R�g��`CD��}�|v]���-���O�(�"�k>�Cr�
�=gzM���P�NT���<�3�l*ƀ!�R��,�c��t)G�)W�����ץ|�f�C����4���pό(q����8��\�wZ���4��sF����p���gf�R7�M���>�s�AE�a-�q�������D���Ueړ���~zJad ����W"�`�,��+ ����T��l��i7VJ��?��:��Yn�( �S�0�k�K�os�}�\;7&'�=�:��:��6�����
F��3�
��QG�{</=9���'�c!.!֕Os���h��M��p�E������ԥ����!���jS?�LG�@���;���,�a9\��M�Ç�'Zp;�g[�z��I��q8���E�� �qXb�K�/��<$�\<���֖$��¸J����+�:�G�k�N)qS
�秃(���8�͐˭gX�\��GC&`C���8��S�Q��F�1�A���8�;,VW�4�]=4絺^.&�8��X�樏��Wk��{e����΄����=xA|���������QtT�A����ʊ�����Jh�X���kv��{����'�i��c�H�'���9 ��,��3��¶<LNJ��Z����}�O�B��j������F�1��͠n"{V�V��y�?N�j��1ï��UT��>�ꘗ���i���k�л��āI��6��+D]Rn����%X1���%*���qcIa��6i��� #u[�F���$d�g�(.f�$�����@
K��'�O#�	����v2�GO꽯��7UoC�������ߌ���X~7��憨5�Y�2)�&�4P
�VM$~�b�`HB�:%j(c$��k����xbqU�&�q���N�}ԝ|��.�;�e6u�~���`��?[K�x?>:H�*�Z5�M~z�3
�q�u}�f�wn���2�sh�D��D���?c1{�}����D�=H0�]�%���]Z���ᴃ�c��"�	B�=�b�?�'�ž>ݚ>q��IK~�������M�1�B!�������[�]��m��lf<؞<H�N{ZX��x
B��t1�dD2�\�7��7��$2�� ê���E��!dlr�����)G#c�(4-���8=wh��$�B��6�}�b�{�S��oh��x\8��
htd��n�su�W0�b�U<���/�? uk��r�vR"
\�7�u����˝+>6Tk�P�� z)����ӯR��"i�(��V�S�"���f�k1���p%���������]��l���Y9�j/�U�_m��Sa�eqH��ث���d' ?�)/��a�����f�(�N��Ћe�!D�哊4���u� NrYefX�%N����I8�*��k����/�6D�Md�̟��.�n��Mp��8�>���4`����p�r?gY4���Z�V����^��p;���tDb�ͤw�׮ۊ. h�EW��I���7��Bs�:�d��}'�W�Ќ��2k)�����`��Ǻ��x@L��/L����X�"@as.��õNj�6�;͖����t��s��?����眰&��&p��̄:}���,3��Ӡ�<��[��
�T�{�u�ZQ]}�V���J��� T�:� ��]�:�q��%܆Fr��_�����:ϋ�)��4��_�{���(��Š�y}̟@���v�V	��LA��!�H����P�M)0��H*�d�9֩��S'���Ki] � dCV��"AjK�G���ʚ�GZ�s�e8��H~ZDO�P3^�݅�
>�Bs�Q��O�'���ѳ��;w�ąLЪ+�\�P�?��
�����a�)��������ɷH�Q6�ZL���n��T���d/��}���u0��k!Vw{nx�'�$�(ܳf��y\`�(���#sÅ��::C���/}ahHw�9u����!p�ehs��=�_������$��7H�|
�s��ya�W �&}�M!���]�L�qȿE�b:a:i�G�x5X�w����H����Γ���r���p���ǈ�V���0D:�ͻ�jvw	��X�W[�Z4�O�擾����N���U�e�w�cW1�pk�3���4�M4Ņ4�:&��ƛXAl�lHL{IX�[��1 ��Z��µ&}��a�<���^�C��p�#Ϩ��}�Iu�˕J<���)��'���Q�(�+6�4��#<Bx�`�|Dpld�&�i����I�]7}�V��}�@��xA�_ӳ�>�+�m�l�2T#ny�6������f�;௛�"~I�%���� �[���S��aqhh��K�!41�^-���d�ŉ+��>�5�����q�a�0�R ���f�z���ƹ�NW�<���p��	�{i��<�6��s0�3����CG~w��^���N�k�0��K�>��z��#�ں=�A|����d	��@+�����vd経��j$۶��ESd���ZI�g��7��:学>J�_a�zp)�'ڱ�T�T{-J8��X._���UD�]���ʿu�i��Z��Ia~O��E�?�\F�Lr����޶�d�67�^f�y�Z�ܶ2�����}:/�\7�[':::4�� g���p�9ﰁ��o���Jp9'Q��?���Ԧh�'#�ku��j?\�s��^α4�Y�Fv��9�4'�� =/s�9�w�z�Em���}  P�
3�'4�\���r�	19,��/0X�ʁ,g{ReNrV��%6)~ءG$�8G+������rY��$."HJ��E�+����py��ߊzQK�A�6#��@7���,�F�,���R���վǇ����[փ�je,�=���z���87�(�I�T�������A��̍�0�,�J��_5�	��Y�ݧ~"9匘���0�Z[fs������a�$+��[LІF��/(��i�E�ǝ�kymZ�i�Fl���7k~��@�w�+���9��x�utt�õ��w��+E�u���x���<��X���#�|}q"���E ����g��%זTYj�I�wS�?�2X����U�*˺o�6`����[�lIX(�fOl�ÄE�� �,���7h9E96e޳pǜW�M�ө�KOD-b�%y2�MF�
��)��
�����Or�R���J�vu��A��f��)�/�3Լ[Ϯ�W��@W����S�5�ȱ��$F�i��C��&´hG��%�6ȂP�S�z6���D��`��*�-��-�o�c_Ӯ�M˛X����g�cW�R�Y!��`��{\U�2ȁ�c�!=/{`e��_�MŇ����P%�WN�P=��Y!�˅:�Q��
*9���k������#�8ǜ�$B$̝ &g�s6�%jq�i���WBب%u����A�Q�I�Ǜt��f*A��o�E��xy�bM�:o�kx5�;>�* �/�_�|i�ܹ��ZC�X���<þ��[I�C˵��@���.�F�5Q�#ݼ���>`@���EA�g���y�}�solXm����FJ���js"�Ε�P;�E͑\Ϧu�L�]��u�A��L�-�̇7癡_{[���������H1�V�]�k����Rs�g���8���m��GR��A�x���-3��\?��XK4ti{���]o���'�IkI�c&��?f��IL�����^+�8ތ��c~5&�4�Gl�%�ǃX��[9Xzh6�gd���%��j�/(���1��+�A4�թ`E�@�	-W֜S`��� s䄿~�B����+T�]��y��"�c�aR?dQ� ,��)�:Ơ!�Ѵ�� ��,�)6�}�{H��2nje��~o=�W_�Nj��׈ti�e��A3��%s�<��G
!T�{ŏ����hd��Y=0A�P�� 3������%^Odl!J/Ϝ6	���L��Ac%��
�&$Σ� �|4D&���հYZZ�/���@� :3�D���]���޿���I�������=%����G%���Kz?/���E��$�eKE]>*o���OH�A �8�t�IX��e�ʖYe������A��F^ꇻ�_���6��@����E�=v�λU��Yޓ�	�[3�Q�q��$�Q���3����lBA����J��ׄlON/cq�\��@�2�0p�S����y�> y!�Hu��q�������������U�,˅����T?�Z�	�� ��Z�ɡAߓ4
�{N�7��=�q��i<��r=�G�Xi,_u)ι�x�/�6�]~A�ē��!4��F�A1�Ft�r� KFc��Ɣ�Hܵ!+�b���/)��3{��K��6�L�s%��R"%]�GJ�y_��������_�(�sW�q��u�c�� ��3�v��B�E�m�n���`-��
�;+`����d"��fQ���9YcL�ĽF���^-G��U����B_�����h�;�Y����0�*�����b{S_��S�z�3j/���A�,4��ϕ��REƆ�ꤤ��j���w/�����ǩ�Q��
͈��*;T��J�Q�b��]˔����+@��f�par���Pr�Z���f?I�Nϔ��$p`�ދ���F>��⤍���q���2���ϟ/�np�DfŰ�3�M�I��B���/��v���v�Q���R޲�i�`�}�S�	�K	zC����[+#`��y�j�$A�*�ưn+G44�:�@~zzz>�f�Hi~�{Ǚ%�!Tz/v�i�I!�o%���<���ķ�����5F�n~uh*�6S)�]��_Uʂ\ԅA��ĕ�.��V���@*��G���I�w���/Lb����9��9��������y/�:ti�sV	��mQK.4!��A�),�ִx�[�msy�Q�7B��?rz���>>7G���ؑ���xn��B�Ecw.�d�${�*�ڍiW�^V�KU��Ta��r�E&)��p9ʲa��K	���x��-�L��@Xls0,���V�����"�湤�ԁL+�)w���q���t"(���2�ȋ�ܥ�Zy�ݦ.�*PS�Y�{E0�G�@���y�)��4�`����iB�ɜhS����)�������/�捉ؠ�/	7=�huPpJ�+rM�z�[ЛC�j��'��l+"IT���w�'�-�W�-���eT�����[AQ�#+~�u���7w��+oX;��*�2L±�Ɵwu �ް`a�n��`�Q1��j�v���w�����tS���%�����aq��aS[�wv�N��4|����r��%W�7��X�R��,���-��@w��;|��b��ҡ���b�B�E���b�K&��y7AFs�~������77&_��zu�mrqb����;�wi�r�e1N�3a���I���\�5@"�!��QW�"	�=]X7r�9�|�����,|��A� ��p��33������<'�M�t�W�*�t�:X d��E�q������+�n���� 2����^Y0~Ju����?��/l���Y�ƥ�l�G��d��.uTV��*K�.;�}��p�&���[vk��&��ps%����z�?��ٹ%h�ݣywN:<�N��h������ia�/��A��ỳ�Z:UTT�p�"���f�n4�F���e��!_�KC	T�c�N���"��>��1�R.� ���T+^�:y�/H|lKtP��?H9��d{��:2%^�3z��z�%o�#���ZG��W�&����d����/�Sj��bZr�p�S�ؾ�0:)��� ��{ҙt�6x��<�=�]c*ĥTB �n�������t��]�8y �����qe�A��7�LP�	���P��zql$\� @���חY8)|����Ȁ|Q�C{��G��e���� Gr�y;PP���߮]�l"���Z�b��}~'��d/�%k���܂�wj��m,�钸���sޙ�D�2t�;�K8��/���Y���Tze �b0���+� �Ϡ�=����C���KEv�����x�a��Kŉ��0��ǱF��?���F�<3���2R�_Ah�BA;y����+���?ի��F-�2�!�Ï��f��Uܤ��/>� U�{QT�ܡ�qdٝK/9�U�3�
V�N��ɥ�7�y�c=��0"�?����C#9����ӄ��n�	��>?����2��N9Ed��?�X��(���ѐ79��F��IFӋ�ȦN��JU��Þ3��E9O����"�;-)q�}R�x�ʭ���m?�t&�̷êO0��כ>ɿ�<������تb������� ~)wD�2�1&W������9~�{_2�Z�@z.W+��3v̌�U,��[�c�tX�j/��w���.K����ҳ'��b��p	���Hd�F���9���@�z�Y9c	�����V\�$<۠k+�k6�sAFv\����������C��t����q܋-
<$Of� �1�ڴ*�u��V�������߈�r�{%��O��%�7/%	`T��9|����+��G�
ı��SsQoph�T��5>x�Eo��Yԡ� 2Mpf�X^��� e^�А�K-�È��D4�B��_l=Gz�t�����~���ʿ���U<�t	��tԎ�F*���C<�ŵAd�N��S&!1CW��x�G�wF���0������cP?6.��Ǖ�[����p�7��ޚ��&���Nm�)x���
�j\vΖ��ݙ��C.D 7B$�8C�^+�Vi�>EbH�f�[oYZ�V�#�L���s����W�����إfg�xo/ZIi)�T�cݛ�o��cB<YtCZr֣��'7�k@Q�g��Ѫ1� ��Ԃ�h��8L�U?�@�8?Ĭ�)��㆏R��5etB��<��M�^��cfj5�z�N�ww���ju�qR�0LS�P|���A�!�x��n�2��=�(p]�_?���=����4�)�t�l�$�u������{o9i�cU�:uV���Ŧ���.\7� v��ٸ�XP�)���lH��ޜ�����y��Z{_G�X�5�:(�Ғ��S����}@�̶�ٚл�1*p�ճ64A�0���B�"S:�s{+�t؛SkDk�@:�j���4���l)�4c���a8dXޟ��<���سŽ�~��G�vw��M<�I��eiw`w��(31(9s
����s����(������XѾቃ��l{��Rn�\/RG�Yc�[ϐ����n���\澴4�ޓ���LRx˱���F��,�u���U>:���|!H���?�.躽T���EѰ���"f�L�n�C�,-FU��O��n����^r*�pL��7�@T�<2�>3՞u�	�ج�wZwgm�&��]7�v��3�y%����7��X1��rNm*��լ����M�KMD�t�0��}�+���$.�z��P.Wu%� qzɲ>��m�R�c��Н����~��മb�a�i�݌c�.�y6;���-*!�A֦C�g_��p��@����4��8�z3���V+�[n�������h��Rm��`!�Z
���.$�W�[T��Mr��/w�*G �gF�4ۈ��8jJۓ���\nPݥ�rMQ��+>5��wڵ��v��R�>m[�Vf���h��w�'_�����{�y^�<���������$�k�~_��;�mt��>��H��H��e��?��SP����Xw�R8�PЫ�~�Lg��}B�C7#8�M���U�b���V�¬i��D�B�{i�4:uP���Uׂ���R��<�J"���/���E��a6��f��#A��(鱐%MH��Ĭ�E��ó?ۮ�*9�P��կ\:ux+s�C�X���T�W`;��sN��'�R q��hv�1��8�~Dd��q?*���Ӎ5��j�+�4Ҵ�"/-2�F�X�5�)c�X�S0�
/�i�g�=s�*A��V���zNj~��.а�E�[�~���ܦ��޲@^��\=����u�cqS�����x����,c��q�;C|�!�-f�N8QbDy+���h|�I�}e��=#�)?�"Y��v�@�ʓ��'/�E�|�Ghʏ�+v�dM����$���Z�C�m���X߂H�";]��j�����ȝ��.��&�;��O9�W�Lۅ(�vK���l|�0܎#���g]dE(ɕq�&�̶��-�6[��`��3��;��2�g��&U�&qSBg���r��;��m�9��;��8O�aP�C?;�`���+�-�zӬ+[��!qI�8)��s3k+��7T�WWV�)��+������4�[��7�]��6�o�J:-�N���@��,�M��UѱnI��]��P���g�cx���=�K�=��E���E� �m��%����"��8�9��kf�+������֓�;���?�L 
8�ŕ�҅��V�H�����H�����e�܉L3���T R��Gl9;*�@�����ĩ2����"��A8`�eH��0�oE��|� �|�H�E��S�MjK�7��d��P>/ ^��:WN�K���������Iim=�&��Z�(�qt�In�ڕ"F�m6�Ra/9�����͚d�]{{���`��v�}PIB+���[#��4[��A�EZ�U�A��!����>^v�W����lې���!����s���G�ru��N=��>T;�m=����K
U?�J�0��-�HLyG'�,�.�F�5{�]b�o]!�(��%�v(�e7�W�W�����5>�͔WN[�����R�&��:_{����TǍ~�7LUL�, ���������֡���|"H��j5��R��m�:e{-�c���P�%9w�y"�:)M��ra��U&�PO`��\��^4�[g�O���ȼ�����C�ɹ�Y}B�'��ƦI��ձX���õ��q�7����l�����	�? �j8?Ĕ<�{X�q�\:Y8HR������� Y&�i�N�̅��p�8��/@�&)p���V\C&�Cdl�wM� �V���I`:7A�-*��1�����aM~�� �"H"%-- �0P�S@iҍ��(	�����56�cҌn�F����|��ϵ����y����_��<�9g��n۠ϛy���G�M����j�ӇY���R>�����u�z� 7.� �[�z�9�� �L}â^<�}�޷*�g�l=�Cdu_�F�E	��4�]{# ]L��/�
2�D�-�e5��l���x�g�JzN���V.%�T���5�G|9�� �%�#� �fI��yxe��{�����~�����Mءl���������_��|�N�;��^s�WI��(�[��ģ���շ��*� \;�|�v�?9��1J�f�s�?K�8`�ĢMZJ�򬨣���B���f:��w��ּ��o��~��{�ڟ�g�A�ݼKݛ�?:��z�۶VS7�`��sj��8U�邒.^�H��(xq�V�@yyz�m�-�I)�A,ǈ��
vA�>������[;Rj��/��鍫�x���7��'I�Y���1��˂e4�yPږ�v���a�����{���i9-\�J��n'�{�����.��˷��	4�ˠ�HJ�=Xc�%��ɭ��m��ݍ6S�Ԛ(�~�O��������u�(��x��S��}���3LDݳ��p!�*�;+��	�N�u/+t��'��&~-�Kɽ�GZC�p��E��	���	h�)��1c�:�u�:I(#sz�<�M���x���Fz$��2f�>���G���X.��� h�/d�#ZT�l+�;�22y�I�'�Cd�m�g����{E�|��=nq����z��ѫ��mC�HD���;L:/�` _�n�*�9XÂM!ȅq��0�ĐK�t�=8�\)�ޓ���?���J�}�@��˱ǖ����5��h�,:���럒}s����u$�u��}]��摵�`Q#�ȓg*��ۛ�*%�������Z�!G9����� ��D�I�@��NLB������C������z����-�0iǈ�4�g//��Z�?LEz���
9��#��'��a��7��L�5ng�_{uC���ւ�[C��W�i/.O��=���(��J�h��Oz�H;�3,��NE|�Mi�d\�;��~�:/�5��	�E=�.-P[`9qN�W �8=n>prT�ϸ�:�����9��W��o	y��Y�t�qT��߂�V���0R��Xn!���ָR�B���r�.Jw��^�gcI l�N�4#>}=e��r��k���:4���W�0>�^p͡D�3�Ӑ�'!:\�XbkŻzjh��G7����,�E9��ID~�,�=/{�A6U�����7{cz����0 ���¡�,@R)q���\U>Jl|�����I~s�-s'8*�;n�n_�s�}U��ѳnc�w�r�ҵ.�<�$Ty�x[�o�} Sg&b7L\��dXp��.���
�i���]U�?e3���oC
��% a�<+5�j/r�O�=�2���ѥ�yr�}��%����&
����MY:T9��n��T��d��og��Q�5�6�W̌ח5���M�*�OB���]V}m�LE�B�����Q�L^���j⋼9l��Y�Pwe?U���I��f�4|��5����WeJ���l2e��I3�g�z0��r��^K.E�������q
Ċ^DR}�M��܂�Yk�%�_��uKىrQ)����[Q�B�q���Ie����/x�{$�t��z�az^R��E[!9�������y�a	݇�{��E����a�Z\���Ř����k߿��?�v�ͻmd�=�}���n$'��S�T��դz���Z������
���E{&�>%j�g����������o-@�R��j\�HJ	�:�I�qљ�S���QҖ�!/��ǥ�T��S��Ý+�L���1�}�����3��n���kF��[�g��������D/��-DD��)�{F*�e��=�%����7l�8�*�HY(yj�1�$igw�sZq�0_���3 4� ���ο�������8��h��P��6��H	�H�[br��7�����N~G9	�-N+^ H�8�����1D�l��D����X���囈Юo���Ogr*�ˣ�e*i�M��o�sC)ԧb�]��C-�m �%�Y�z�fD�g���3�����K��^���=Vs�"����\��u��1��}9c/�[��N�z��X�?�eF���]�nF��>�UkY4�9�gψ�ˈ�YV�����ڸ݋t�ͷlI���}J���gMM�8���.�|x?��Y�힟���k�憊U�qC���A$��ϰGֳ= �e�+��i��ހJ�2,��ac�ޖ� ��ė������'�=��_{HJ˶߇x�o<���U�|B��y���j,���ݲ�`�T��H(�n8�V�&[qdx�S��\|��s����w�G�-��ϮL�yx�y�d	�%�w���s�)tzo�H��͹?���6���F�[�$$~,�~̴� 
�.��Tj�n�,���`�ѲZ�7��"�CO�:f$�����D�����-���d�����'��⧎���m�i=a*}T���o��'�L�	����w�0c�rRN?)���b�G)�&���3�]�3��,���9yZ$�����KjU�a�w���t22�V��F2����l�9_�{�͠�i�J"d,[(i��YfS_d�N�sui�̬��^κșs�}��SPa5-p ^�I�s�[9�C㭶P�數zvw�����=�l0�{�0�KCbr�l�	�����j��ì��*�(���&��\N��8���� �	��>��L>h��"��RIE�i?�;����6p�gQ2]x�J��N�($�'陙vo�5p��#�
��Q3r�Ch���2�QU��W���vf�:V�����'��/�j;°�e[p�^��P� 7d"���ǲ���sxPis��%�絷���ˍ;ɲTQw���8���^�Ϯ����w�Ҽe�w�-���sw@�?�`̷�ZI��j�i��$���D/4X�FkfW\O̡86�ԬKЄ)
)`�q
�e�B��4�}Ob�e�;|[��G��Յm�aq�g�tPDGb6�05���)U	��.+���!G��5���O�=<B�Y�O�mm�@�Q�ȁ7�����]�z<;	ųLBS�k�$�Ԗ��?x�[�YcF��_Y��o鐜�M��q��څ:Q�J3i��p�~qJ�Y�;���@����K�L�#��S���|�h�����d������F�zA2㊔h�}br &`�������L�����W�x$fL�f��/�ǌ���S���s�%���+ �/�����Xc}k�R��*&���F����z��g����zc?��)��.Dkh��� 8Uj����#^������h���q�-��&���?�,�s�>�o�,xI��e���is��̦""4ݳDz{�H��~te�\rY/#Pݴn�5�>�u[T��+>Y�W�e7'�7REI��H�r�sF�5z�=�ْ��nw�<��<C/�6�Gb��_�e�ܴC�.�[���
4�ɥ�T��]�Y�d����А��0�9PG2	C���̑m���N\̞Ϣ�^���K}��w|�t��U�D�{�M~5��V|$�ɴ���*R�W�Dk�ݚ)�&��<�:n#�����z���B�PS��J��G.��'����x� �=�Pm����x���5.�v�l���l��(�|g1�l���̅�.�.�������L��խ��ݚ2�1,	!��l��!&<³��"_G��k%_�9vN��1��z���.�oc�x)Έ�6ņ����]�}�6,^�8u�~�|���X�e�
cJ}��-_����ߗ�뻗�;�R�[ 2��q��2-���'7[�9	�c3N6e&	�s�i˲��S6�m�!wM�.�aB�Rt�O�R��[T�L�\3��m͇l�����E�n��T�z�2���#�?�3�so��I^��]jFj������¾~�����h9�V˅�n��BHm���F�dn��^!;E1'jkm tR�ߦ�"#�S����zC�@�����ȧ���ֽ���K������m�o�aDYc,�O�؆�G>y�y�L��h�A!�B�0�aFT�eS
F�1GӤ���'U��@/{�<?.��te���8��gJ�Y�s�z���1�l��$�;�QY[��_LN��.� ˖�Z&Gu���:�pR�S��ޅu�犜��'m�ݏ���g�$#���""�b&�/f�$���[�r�f�j<��x) p�d���ϛ�,���S[��"v���9D���χ�,�I�m����R���U��B� P�oF�U�3�}M:[��)2��d�O9Xx掭��� '�t
�����S{� �{L\L)��o�)"`���i?+��z�v���(<6>��ώ��-��B�G�/�^�џV���yTS�Jͷf��T�pU������� ����	o�	�V>x�/�����*#�ڝ5:P'=���]�ݖ�N%߳�#^kA����xT����!��?��-F��r��G���ޖ~��̙�)UX���IV:V����tS��y��\���>L��Z��݋�vgv��H�����9,6FW�U�6�/�v辞�y��ަ��m��/�ʽ�8f��1x)�+f�?쒗i������wy���kJ_��� �3�*��Y���^�z+�]fa�D�\x�?��(�y���������ß���+PϢ��nߞ �̈́�`FJ��ֶ��4*uJR��u��x~踶*�+�~��k�/5��Z�8o���<������k�!�H�N���������E�-��=[c�7t��=�ǝ<���������gW��c�Ԗ���D���Y��G�E�DF���7��Fy"��ワ�%�kL�&�1r"!�f)e��ǋ������co^x�e,��	+�.���sI������s��~��E�-y�\A	mFM�����M��&�vn�}I�w����r൥�]U���{��.�"R�HO���兔���S��r��&��/m�0�e'y���;�<0�<�I��VW���$F�,��!���^��F͙N|�̶�.���o���s��&�ϙ���M PjH���B;�������cpl���U�;�*�����tfͩjn�U��ڗ@F���{D�AW��#$���o�$F*���Pi9r^�.�=�	/��u?���{��qZ�o�s5_޸�}�fh��#�
yߦ}� ��Nt�Zs]���4�,�u_A�:�hR�'�j8����<��.�c�l 

�¶m�ͥ�T7N [0�cE�GU��UV�ќ����d(~APl�l�Oc79�f�rp~27�����m?p�������z,����sة���xʽ5�n�ߴ��	�2�0��砽�(��ʐ-�V�� ����޽`b��;�])�z~drhh(cWW���K[��k�'�p���g��;n[�N�w0� �'UpO�����ĕ��W���d��^f�Iwn���+������ey�����z
��w�n^�bK�r�s�"���W�B��x�'}Rٳ�&��/�(�}��t'���4)���Qg)ה�P�ѷ&��������Y��Qzڨ�ٿ����j�O/xy��Q܈��(�Y0��ݠݚqW�y�j4R��6_��2-���3v �9;{C��|ܯx˙��������{Ny��x��6&��:5�A�;�w��?o�lu�V�Rb����P�����M�Gwg���:�r��u�fy���S5Dh�J��E�m����o 1 %󺙏�h�G/)m�l���#�]f�<4���[�G
�Q�ڑrMe��<FNe���Ĝnx�>��^{�d,wz���W���UĘE{����f�7�߯d2)�4�����Uv�Q��h�1E<�a����W�	�[~Y�=L1�}m:WB�H=�+��%#�ss�S�)w���[����m}�<yl����`��[ie&�0O}Uzq@w�f�SCWdсc1�k��*b3�n�S[
�^��P�Rz�Jfǲ&".�Tȷ�Y�B]��f�f�Q�,�bhRM��o䋙ἤ_��n�o =!�R ����MAb�
$��0r����? 9����<Cwg�+7+�2ԥ�GɵF�׾Yvηb��#�Ut���dk%*?;��k2i���JE��d�=����S�[�\�v�;c��N�%/��V\,<�Ҳ��< �߾�m����2�ڶ�Z���kɐ�^&ܬ8��]~hχMXG�hL���W��ߩ�@xZ������Ϟ�����Px������BKR$�U@�~/�`]��Û�$e9b`����d�25e�&�L
Ƃ�Xh�����3�_(P���u��,_%�d���i'�M�k��RP��:��DS�����툰Pb����ßO�8�iv�䃻��M>_$*��5�_)͍9	NW{W�[iox�G�7KEZ��=ܡCo�
2H�����ޜ 0x/�tϯd��(1:������d+(�A��f�e��
x����L��m�ܳy��D���������0P?wn:<��c�r�Sc�.lr��=]�.b�M���Mϻ3""`%�>"p�&�f�F��nR�<�k����*V��ms���>��\L�ܑ6�n��p�gR��*�G|K�aJ�����;X�}���K��#���M��<gY:h��v�2%Z�T�#vgE��٭��k �t:��;�_䖑g�4�9:�����n��q�C�U�v�;X֬�!:��r��JD�~�l6K����kF��V�^u����T��B��F,Ssh�3�-�YT����/~��ސ��"m�=���w�a�ڣ֬��Yc�Z>�� ��}�r0��L������J^���)C)�s�_�r��Զ��p'1QX%�!��)QR�2�Fޫ�E��Z��$b�1��W�t�E.�"��=�(��[o���@ �%�p�a]E��̫l�m]��I�T��]����O�Sx]d [��x�b�>�JP�"��h��tP?���1Ҧ��lE^��(����o5*�~�&���w�m��m��0)�E\1�}$K��C��#(u����J����gd)��;p~�t
ٹV>|�#�����=g��$0�,��#l�z?�㒝�նb�������(Sz׻�'�����˂r�\/����LH�0�����=9��]�aO�/��tn�J6|O�׳�"`C���KF-��M��|e����5��]��	������1?�]qD��iTu����S���?��@%<���x�m�%~�bB���-��Z*��	��^�s�د�f���m�m7���=Y|���h�׵I�4�7�ѥE�H��aR��f�*$b�������Nv�-��3y�`S�AD���/i#��S�����\��w�3E�pj
����Qæ}y��NN��d���Zz�~��ސ�߼�wې'�j{cV-F�c�O�mX��o6�?iw���k�:P@#��d��1��۴�
�m�x�>$J�-�Z^52S�ߵf�-�P�ճ��D����������cUx�6�k�K�+/�t�d��W�:�^':�{�j6�>���v2�;�x:��
DԪ}.�M�y�@�:�QQ�����Vtmv�w�e���л��}�=�5��R�����9dS�������IEj�d?p��w�=�cQ#���gW�k�4�;���[��ƽ�%E�or�[�k�K[�.&����{��ҵ�H{���������ly2�k�(dv���	JKC�����]j�k,ң��պ���X�,�hH���������̓�mz'�t㹮=�`k�����|:N�|r>�C����7 %3�z����{�QT��T��w�O[W� �ڰ������R=����(9���§�M�DK(a��h�qZ�A�����	@hL����vd���Vћ�ƛ&b�0����>��'zbh�K(���s���Et�m"�ɨ��կ�QJ���XsZ�_w��-j�O��'k�e'�ss��ÜQhC��O�'���}D�A�@-|���K���ڸ^�>����	�o<W�n;�7i�|�5�'_3J�>��.`�9����yL��uL�B�{�RlB�s$�@b+����NNZ�� 2db�qJ쀯���ƃ���	� x�+q�>`4�{��ǡ�%m���C��/;8�_�G�]aE^�t��ж����]ܮ��w���������+���#8��P֣�/O�����{��\D6@u�bꕖPmd��q�%�����S�}��)*@�0#G�4:� OQ�:9��ν�b�Z/
i��<f�����!����m�+��Q����}~�)�ci���ޠ�l�Ԁ��!f/�X���"�A������X==[j�`7&�DW�<�4�ֿ�C`ߚ_�錴vi��k��̱��/4Ɨ��^H0 �ҢR8~��Z���"q9gr?4,?>�Z�E��aF.�L� G�ILKo���y3Ju�f9)o�+T�`̊F{�jJ�<|H���C�~jK寂kT�^��<b��}���h�q�^0MrA��<�)����M�@`2����f#�^����¸�$�����$3���:3xZ.}���ͳ�юvM�ƕ.�M-���w+���� d�C��܎�zp�~9Z�e��dR%�E֙5
�D	@9K�eib��｜����'����{e��]-&�R�X�6j8�RƎ��Q����^=M���s��O����"��m�rE���Y�#^pc�h�h��D=Zo���MQ��4��x�A��'o�_>BN�(�:G���0-��߽-�.�뢚_R_�ܝ���z`��9>�Պ����>&U�n�>��(����;�q��-20Pt���x��w9�Z0qN ~��N���u@�7�����Q��<�>��3�f��yHF\w��%Ә(�,o��R,��b�E��)�e �@�5�TB��:ne�B��j`nC��_�q����5�^4��M����GͶ|җ�֧\��'��j�U�2#��%��3�<�;]'O�BL�ڟ�O@+*h�p��II �$�n]9���{�eU.*�O�^9;漬V?K��=�2~��"�����d�RTf1M�����tJ��G�6o����^2D�;��ⷼ���_;u�B�d�s��%D�e� �G�U����t�F����?�˨�'9����΃�S�t���O41���c�<�ڈ�7N
�R����Q�u@S�}��������y���[�:�~�#V
����N�@�lK)f{M�6',p��,_����+�+�ƚ�'G�h���K]�8����(3��j�9�`�_`��ޢ�0�,,�{�<����h2��K�&[}���m����v�s�)���>��?ε,�\Ze�>U{hV.a�B�c~3�� �I����]kXw�Kw4��Z~.�F�t���[���?��ޒ��bC��:_&c1��������M��J�����4&z���^�Geń�x0���\��@0�y�66i�,i��SQ%�r.�子&�p��/o���ר��{G�����s�i���o\�<����\"�˅{Bj,7<�-����h]�B{���C$R�+`>�¶���{ ��8���^��引�K��ׂЭ�ߊ=;"�w��������#���o�d[nu_Qm�Tw����T�*�Z�Y�
F�b��]�l*,�jx����=N<�ѣl��KLQ��SNNR^��<H?}2�UJ�5Y��?�������5��PO<̐}�dS�@g��6��E%���E�q�@��1踠�uFS�	��DϘg����5�r1c|��/;a��1�e�T�x٨�/c[k.��f���U��7b։�3��̏���G�R=���KM�(1�H̺p�b�w͋�����QCn!�d�@O���3h0�x¤�EǠ��&+>�&�Qlr	���Fe���lWa��Lֲ�P��{�>�B\�M��bBrmUD���_����"d�#g�{�q-?Fy���������	�+|D���,�l<�A3q���<���lz����T��X��2~�����f&e��P8Ru8�z7!q+֝M��,�	跼+��gn�^"Ϋ���?�ژm��Z�?��t:,ifp!����`�4�5��A��~�IpRY�߷��j�"��7���������O��;�Ӻ|(L��ė��%���nTS��,CGe'(Pz��)�YK�k���Td媳�ڏ�Y��N������i��wr���~R�ֵ(d0?��_Zs^��9���Y�/uk�q&梁��ż��nv��b�te:�7/�NH��a-l���sssOn��D�`U�8�/M�
1��S���;��#sqE��m��8$���M��G�B_}'���~�a�u�8�iq����I�nG-�{��qttR��7׉6��Z��a�_ �,���+8j��K}�8H���'/��O���}äs��sW/�l�O��5˱�݊�2T3�^U�o��,9bD^�j1W7�������@=H<#X����f����=�"Os*�K�'צ����� �����Oacn<���ṅ��,A�����jq���O�wd_�����7�觿X��"VE/��lufOl`b?D�����酡ܞ˶�����e?�?7 �͒���w}_�E3Mv�Ǹ���i�!��_��/��جt�Wԏ�*y�|OЩ\8�D�[�6o��o��'��B�b�_�:����p��B�nBL��Y�/R`;}W쇹��#1�I���_ѷ�7� _��s5����u��x�CT��B7����#���o��0���2ҽn�t����M+�|.ݽ>LL����h������r�����F��gF2As�-�
��Ʊ%���=�۶����+7+�s� ��M� nЖ���Y 5Yx���7���}�%�y,�b�l?�{����L��d��Gc5����=L�b���h��v3O��L�`��)���;��a/8_�y�\R뼵��_j��tk))LJ��i�{�	�>=*�\���غ[�%������-��(�>���pm�s�0�����%x4�7M����z�����b�2'kĚi�3����7����z"���I��#���d,ҋ'�|��5��D�ZZ�u5�� �{���q܍��Qw=o]�F��^�h����B� �}F�1s�c��ToUlK��^"����^�ǩ�������o���^$2��T�[�#����,nZC`��ѣU���mOE"*�9���wd1&V{����%���Q~T]c��8�Mª�('��=���]A��7��H�.-���������JQ��I���M��QM�"q
�no�X:F?�Q����/��{0��=?��-	\�Ab$YM�V	���^oN�'E��7�g�d��}I��f�������:��I��3Zil���S��\���[ 6�>�]��?���Ay.~�����[�*.i�)����>E�sM=�=�"Ke���gzi����j4�<3����$u��AD|�����j.z3 �#��Kg���8�:��d��{v�C�v�mcF��v2�/�0��˾�1�d~4�2�N;�����el���G�Q��c���r��Ͳ���y�$l��_�)ז=�i�~8�5�
��/�� ���ȦcJ�9�T��w�';����e�ͷ�$!ϵ#צ�9�1��KM"�iN7�YZ�a�V3>���U�mݽ;?C��?�x,,����M����3@�r+=(��;��-LSJ�L���#���7�ۑ6i��I!/��>�Gi/�j*�ҿ����bk�F�n����W������g׫yq��?mrA��T����y��P���rCb0����}Er����5t�9�	�:RD�R�@FL
�W���tA��]j`�sO,���]�F)�A/��]#��bDq�w�>��<B�.�cI���Wu��ݘ��x��ȗ�5��� Ts���%~�p.��eޚ���!��0��]N����^�c����\H�b���p�q�g#넍3���?z5����\�^=� 8D;g}/�x�mf�=zWAy��N��~���3Z%d��Q8ǃ��
�ZV��
t��
�����>������a8mp���]E���_	$��B�AM�^g���E&�10���jW������`~$��<IH�6�l�ٶA��{��_#O��?�#�E�F�8���8'���7f]��A�:'��Q��][�g�ƕ���?��nv&���{�^�x�X*�=� |ʟ�<\K�����_sAH-j�|���N�ֻt�yc�f+�XǸ�CH�]�Xw ��fK�yx]qR��G��φU�Oq��SRGj�>���wV�,g�y,[����w��*���ZI�U�`�K<����K�P�vV�9�TM�U}HY��6���7b%��Fq<��pSͬ��gxw����̞!����w�Z�O[�4��|Ѵ~p�����������}��$��5ȿ������h������Z��C�d�6�\3��z�>�O���٨8A�F��U��&�����ѡ`�J]�&�� 4�$���\�N�zoR�UU�	�Z���I�L*}�5"�x�}�Ӷz��1Li_�ќ����7�HD��P Q$�jv��~��j�pV�L�|{���c ���W�I??��T�ۚ��P-���M�=�O���!\���S��ʛQ���s��0�9� d���ydF1����,&)R�ϻ_\������}���_n4/
>���̖H�t'a����<*O�M,�R��ڲ�Q��8��9���ɐI�"�"���v�¢Oh��8!d��w7��H�0�����.NK�����9*5�0c�rb|�pO�D�AV���6�Wd�LD�Mt�
�ӏ����M}��Jd�P�=i�v�R��<�lu�sﻬ$hdN�K}����:�B0%�<>��/��E�UD-ɥ���������8�5�/�D��Hش������v�e{��{�
'b����j�m�9�~H�8}����*�*-��qR�x�3�.�;[7�<�a�~Y�T'd#�ԑ3m�s߶6'��3U��s?�Ts����e^Q���~w4v1k,�f{ Q�$�����ɏWMG��	���jO�����*���h
Op� f���J*�����r�_�W�(%����q ߪ�7�=|�2�Ӂ{c�rD��t4�YdcF�u�O�0P���(�8w��n^|��3)���Z#2'�5J~
�0<֭t�����V�m���mމGzlI�M3���j�@����`1,b���v���(J6��P/,�댄�a���;L%o9[Ju�d@��%�Ȁo�uI�&s_}y�] ���9d���aTU��9ϥT��>0��Id��j�3��^���&K+>�����"r��J�����l��U�F�7N�֡Z���f��Q �G/�j��c_��N����������s�|ا^��cT����"?�<I�Y�E`��cO��!Ů��2���{�J����E����@w��W�N�1#�:!��
҆'�d���bB�M�f���pY�e6�9��#
i���@^M���-��*�Έ�K!`N�VE���/b�8�B�kj�����֨2��#-�����c��\P��O�h1"�g�~�֤�qөP����NI <3>�p�^@ʹ�3��gt4�=�B9-6���7ٮ�
]��)��j�z8�\�hK-�7�jp[�+��z�����:C�N�fEA�ٴ�q���X�����ܿ]��|�W��wc���T�'{��z[���IG�H���uOU�Cެ^?~�;H�X�X�z�*�e/̌$����Ÿ�E�Qv\�2"���V�F��2e��cK�\D�$�Օ����Mz�Z��l�TdW�B�\ū�e�v��כ��$��yLU����9���(��������5q�̓�+.#PKj8m �I����.v����jЧ� V�@���G$�D�����҄H\��	�Z6��9yN-��l^���]�bG�F�B &��O&b�'����L»�e�kU�L7hhHc����sW�����,��-^���j�����h�uF�'}���f���Q�k��l�wgO��W,����I�a���m�3�&tQ=11ڛ���?@����w���V53o�\� e��5lǥ悏�K��i�tde*�N���T��,~���$nb��;�n#Mw�R}��'D!��7��{V4;�2t�*z:,��@j>�D�a�YI��C��짬�c�;�Q]�Z��%CE��g۩&}��Ǜ&���I��eC�֊��.�N3���h�$C�>F?K�F&�����*�����XY?�>3n|���S�~�s#~�<3��fk���|�m��z�[z�J���b9�a+?���$��V$o|An�y�.��^�ힲ���3��;p1�wp?����G����{�L��X�x4N�u��q4�o�?����Gj�}�t�Np[�<@�[����f�'Y�]AS�C���/c�v�HH�����a"�,�5z$��p�7$��K/����a{����[�V��$iR]X�e���읋P¿��,7�ԕ���ʧm��W&�|.�V������*~!����o̫��o�������ם��S������KW�I}���'�s���JgR�s�f�$�Ӿ�^p9�#?���DR�p���g�g����,�,[��݌�XI���h@�1���o�L�->K�dBkO�c5��^>i���YU^nU��ͪ��s_]�
���I�jh ��S3����mV��k���$:U_\λ�A��m2 9>����h�"_f�Z���H�'�����R{���8��'Pc���W�Yz#8���~��e�����8>�,\����ʒ���c;��J[�K����B��b�cE�|p�X�'k�p,��� �ε�27b2���S��^i�P�m�|�}��� D{����~D����}�f��7h�[2Ǻ����o<V)q9dW:E����,�1��XRi����{�ֈ��%]�?365�$.q��p�ߤ'܁�rd���!�<֛q��>M;��&��?/D_�IJ�"��g���{��\�� ^���U.R�_3|K*t�<"�>Y֕tH.Rs��P��3��[�?�V�1P�b�̚�q�@���OzT	��rH籱�R�0��[���Afoo���(�	*IĤg�놉MS�D�o���ǹ5��[��0[8���J�&�hF�f��Og'��E��I�2Tpio���S��}B�{���|����\/N��Ib����C� �S�0�38::��/:a�k��3kTf�fs*y��Ze
����m�],a�Rr��HV:��_��� ?]ز�����\wI��<y��r������)(<�h�7��lK������'_b~J\�V�y��L�8h;C�Dl�o+Q�'�	��Z{j���¢U��jDm'SN�Э�����K^�:&8�$�\��q�w��+ �k b.06s��|��_�B��_5A
Pi��/�	�ޟ�4�z���sΓ�S\�l|X`�#��ŭ�}RX�_(@um~'�:\_��d'0�+�`a=����� �z\~ٯw�"V_�7����ٞ�JÙ�?(��O���A1�s��e���|߯Ƶ�R�uS���$�r/��@f�Ag'�Ep�ì�A�$��d�|�b�q��|�o��Ywbh>ֲ�[=9e=lh=>�`����z����nD����N��D�
@'6Dձ2���-��?���z��Dv짟�\��G`��b)��wD�>����Z#���Y��$���#'1�VŤ�rɝrb�6�[�ԼnUͦ��a^��z�mg�iȻ`�z�գIMBWq�p�xc�N��5-�j�����7��uj���C9m�Ҿ`�)�~�����T�4t��Ħ������#��V��a��tӍ'����~�+%�mҔ�&���FK4�6O`7���Q��"���J��A-�	p6�ϨaO�R��{�`uK��V�,����t�w^�D�UN�����^tܼ�S�۹G�b9��b��Ղ���|�+�K��?+xs���yr�}va��u�+�([	�k;���l8 ���O�I�+J�j���w|D�{ǪF�:��hU2���*�1�LF1*\�I*��$&��l�m�A��;���j	s��/�o���m��~\�ZmXT;�����-��~4��S�Ac$̗�Ay�>�Yr��ˌ�.K���ջ���\���/�x^3����_���њĝ��7_,�Y������ ֭������)߉��Z����z-v�Z�3.Iq�+j�J@d��nhzl���m�C!sX��`hz⌅/!�̮"7[m�K��Ȯ��Ei!��E߸���B����̀b\v�D"�,�WE�l�D��B?�(���;A�.�%8�`ae1����rc_:hHm��0Fˡ�ݐ��uY��5�f�NͿ2T��5c�M0F�^�~�M3�׆�
�,v��3Z��T��׳���EC���,� ��`z��
�O4�.O������7U�k���6��]��&�n�J����JM_�ϝ�i����6�wm�t}��^�y���>�,n��ɯy�;7���_�9����ɏ�u[��޽o}��)C�	��(p��|�d��`���34�����`���_N����o�������)�	 PK   J�Xh`Pҷ!  �!  /   images/4b60cb4e-ac73-4aba-afdc-1cf5937e57a1.png�!MމPNG

   IHDR   d   o   %e�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  !?IDATx��}	��u�WK���hF�h4Z@�b��-˖B�b�����!���'�|b�CVs�3�q�#�lr�y/��`�1D�%����/�e$�F��=�VU�������Qk�A�{��U�]]]}����:.�<��c���7��;�a,�4�֭å��>M����O�Υ��KHQ�O���3)2�d��<���*g��{��y�>��2� 1-�C,χI�!z�����P	"�?RTbA��C��Œ��_�I��T�j<��0z�J�W72� ��O�Ua=QQ4?,����,�2>m!6��+����I�Z�U�����˲�	����?H��������'��@�jڿ9>�Ĵ��ʊQ*KFS��ea,�z������S<��2@!:�
j�Ytʍ�sc�O6wT�8҈�=�����{��8��w�}�V�2b�ب�L�"룐�,T�D0sb��zz�a(��.�sF���0�O(�	����a*k�p˵;K��_�#m�p����%�>Ҍ����6l؀]�v�RK.@�	���^ȅ�{�8_g֬Y�����&�Ju,�����'�Pۉp Ο�Ce^�Ч�9O�8?����ޡ�q��Ӓ�Qۅu��8':k��D=v7kN!P�J%C�6mb�e/HL*���7sRKe3��Y'��(�?�>�����T,���� �($S��,G���0�
Ź�|O�f d	'�?�"��_Ob�V*g0�&��Ϝ�_���p���~\<a��P��J���\��s���`�ԩ�6m��p���25�J������J�ta��J2��aZi�[� �<����{��r���`���l�[6`F��d_��-i
��G��3O�dP�rr�0u�g�����#�����CKKr�V������{0g��~��={6�� 
_��לƲ�0�B�Gɘ� +c#�nҫ)�Qt
�BTL�Bl��^�}w���ߢ�M
��(����AX����F��Ə���?�#Y�h���_<����
��u�~l!NuO��-r�*ʭepp[�n��/��H$�Wǎ�թ�\�w�u�~?���Ĩs;�r|E����� ���̙x�n������R�H��5�� z��T*����X���<��f����z��o�rV�L7ӛpk`�4f2��P+�4���F�{t��%е�[���R�r�-hjj�������9��c�p�B�}��B��d2�3UU��x
�3EX���gnGyh�H�@��l�@״��9L��_5|5���~J7��`
,�m*�<F��p R���6Q�lW���?��0�e����V� �\C�]�C����e��?0Ps����lm^�#�3�A�Ȍ��c}���=�Hs����җ��G}###�����g?�Ypu��X�-���"�=p� ��������9S���g�٧$P)�l��L`%h�P��f	��T� +.ML�moJ�+���
������
v��?1o
���*�����9���>2sC��� Fq(��"��`km���N|��8�<��OÄ́	¼744�֫7�,��������/�; s��E}}}�E�)�[o�%.굉�����+pݜb�b�޴�����B�@+[Fe1_�� H�l`V �L@<L��Ҧ*�Ӡc`J`$8��a�#̚9���yG�4b�e��B?kH������5}��ս8֚ru4�|�0Ϙ1#�����+��k�axx�� a����ǜ �������wމISf ��:�rS'����]aY�c�����V~��	f�6	�������	n��l�ထ�6n����[���SP�����ί�gYqGl��aa�Pp��Z���F���}������w�^9r_���l�2����"R=x��R^^�q��Lm޼Y����_��{()�ƒ�q��(���Ri��[�Į�EЫ>*�QP�M�'�$s bf1$�\yؑa�4 �!�4;0��B������S�V}3���`��F��(���n��=�u���������ß����o|����׾�5a���M?��$/ �E�>�o/����֮�]�E�<�:��ZrH�"����K(X�M�^�Zx��"&��4� �ad\�F�������L���$`�ۄ�?���V�y(%Ka���n�s��(ߒ�?�'�o6��܇��	qW�x��c�쫈$T޷��$P ^vp4�g����R��@	V\}�S�b�*�L  iE�G�j>N/)�����61�$lP���<�ʹ�N.S�M�O��bbQd���(A�p�!��撏�
�ޗ�;|-Ä�(�������W��+�濵�[innơC��`��Q��9�-M��ٳ�[c�e`�h�Y��#���]�l�"�$����$lF\�ZV��0�I�[�,v�6�
�P�;�c:b˄����F�X��Ӡ(�������Cs���>i�l�H!
�� 1===b��;j����H&R�1%6 �(���u��SE�D�C¦��5b���������c
�i�d���d�b�1%%�c>	$��F��$��$"1�|O.P�ML�H�Ϡ��M�)V�p$��][����,�%S�� B$x%t����M��`�hE�#��φs3�x��J� �k�!��}���|Zd�x@������yhi��h[4��%�1�����,A�����gP��Pb�x���iX�������b��lSŬP<@(�o��EJD�
�D���1%��S�����gkºoi�J���p�����?+�Ԫ��do�j`2�q39o�3�n��	0"H��'0�b��
��*%�!v��43k�d����
=��!|�/k���I���)g�km���S+ېH���H�+�uSX�x=���]��~�6+>LbH��a�l�v ղ�!@�����]"[[�O�X���nJvc�!n���n�h�9�����F$�D�3o�2���5Č�t�F�]	���e�Xb�1�aa�C���5�UQ�rE��e����>E�f�T,�~m�q�昿�?�+���3�7ǦK�`�[�������D��:�W�a�>�`xDT~r������}'+2��$�͗Б�8f�Xn?Yq�{xu�d��|�no^\���rP�(0�T�kn������}<�z1m�a�
Q�#�|��TBWC����K���KM��**K���q���'y�-k�܉�o���p��ĵ�Y��"3������v�n�d�`f�0CVj��+�u��N�VةϝvS�eN'����ἀ�^t��V:�s��8\/E�z�"�u��%o�ʦ^�������N�ZD`��NW/Y������k��`�	�����B�Ǎ��D�j	92r≎+ ��d3���긏���t}F�3�J�M6]
���	��:����͹. �����q��3�����
	3�`�A���zi��Ӷ���f��n��t��k��wh��U��~��e~�Su���/�>��z��,���F�N�5ı�wlv�0m�A�T͓ܠ\c�e��X�M�e��d��U�j�Xr3R�fȶ�e	W�/�[V�j^͉ɫ5��}{9��d�SU�,�(��`G�+���Xr�{9���-���v�_���ӧA-�V�<
��U�����z�M�q�&h��K@�@\�QU�����f�.�h�꒶���Z���ŗ	
}��fd�H�-EqYb�Ĥke�b�zI *�@t�M�% �t���3E쨧��O�߸��pDTLF= 8-����Ǔ]���?�2�%�m��R٩��Ldd�b	��T �!.�&�c��R���2�"�F>q*%=� b���b_-����.��Xܜ�:zز����5�-�"���z�\١.�z����4ؙ��a��M%&� 9[ٿL	L�2����Y<u�<Ҁ��m�t��<S��qkq�� 1�WZ��zYU�\D����.D �N�oM�܍����x�E�= �C�a�j��U��r}e�Z z0d�zE0r����L�^4	�5t��N��v�39�K�+Ki[/MT�ws��N[@��"�[P�r_��$��}���i��fk)���e�V�[_�1[z�NG���%f&+�N�1RĒy���]+�֨���J0 %�d�ntLUڡ�b܅.ƃ|Н>,����O�أp�{�;����֍��hZ%��&i��+S�+-��CG�ME%�Q���ȮG
��W+ǧ�f��IT�R'��$�O��?�&Z�_�宴/J������so�@=a�"���r�-�=k&��&��*'��}-BQ�Q���Ng����������&����M�윬����E��o�q�x^�	�v뙛&f�ˎ�҉����~����f���^aw��s=�WH�0 ����'�R5���8/�e� �C�����J)�)v:;�Ap=��:˭PLGY<|@!("r�"L~*{���sv��ny*~���:fHE��t��\�Q���S�4�>�BQCp+u3���H
M�!��" �.�3/��$d�D�{Ve-��!>'ʂ7�R�""�N3F��(9:�Hl|��e�����${԰�!��NH4ݮ'Q�]uR������[r��-�)��[i �¢�����d�i��+�t13�i�]��t�1�("r1īC�)s�In�2C��T8��a��LCދ"J�p	Q w��O��MgLKw�v ��&\թw)�y�[5bOn�U(Fy ��(�4��$]m"���b�Ʌ���cTF��V6YG�]~�͸f*#����""�.9Ə���Ԡ=(˔I9�N����{C^˰���WVS����;m��G(��*�<-�(��p#�]H��kY�#(6Q��(�TQb6���D<Rw�.��I�~v�9v����kKrx�����h=d�\A�423u�"\�۬G{���fQ�Q>���~$X��I���p&P��C�g�H�F<ڮJ����)�#J�o�$���L����R�(p��r��m���z���l=�v�El�ퟏ�.���p��;G�=������&�趙�F��mU��tB|��r�����Va‡�`��<f���Y2����&�ɹ����u[�ܜq]�#�${��\4[��|�L����X�yݖX'M���V¡��Z���~����>�v�J@�R�hȜ�QN#hDx�~���S.K~�$��OF��H�{/���ȏ�!h����S��@1u�3�i�L>E�#�H�ά��WH���9Ч��~"�����T>��<�D2���S(��T4[c�b�"wRM����vtH��~%�[�D��Uo����idɒh�I�Lj��Y�ODt��6L�o��N�9��?��^"�_P�MeQ��s�a��J��-�$��&J2��j́�b
s�MXv��ZQ��8fKSya<A��{fvu}?�~��z2��"KF�*A@��"�%s���f�)�5���<�� ]���/�IC~�	8r/?p�&T����0���:݌��K�,���ò(a���-bG?��(��RAgOr��gZ_�;3��n��^��Yb��H!�����3Y�I��Єi�O���+�`w@��y�x;�c�Xa�a��x��*�����cO�
��k�+�\�����8���������I[��f�Gd�S4]҉3j�`���y�������|*v��w�m2���Q��#q��C�x�~$��^�aH�c��0��M��j�H�o����R�x#*Q	����"5���YVh ��ޖ��I5�o`d;x��p[3���&]٦K)I��WÌ� [��O�	��J���h뙆�-ܦ~l,�'�$��d-n$F�ⲥ8��4}Z�9�~Y�%#*^9N��U��H �M�^������X�-�`�ѥt|4�U���R3p(�i,,ya4K�ܤ��T�[q��[R��
�V�$��EU}v��qŶT&�=�]C5bպ|2�Dʼj���M����$����+>؇���jε�rƓ�����`�$�I��X�:3#���dO=���GN}l�>& <~��SvG�A��P�r��>U�%�+Ἣ�t�M��
��>Y���~���T6�ALۮ�e5���Φkؚ�'�k�_�<���#?�t�`T4.��Ay1�c3R��3|r)#�/$;4ME4����CCMC��8�5���-W�+)<�J/ΐ/z��L%G�[��~Bt?�d���2s���3z�0W�nf�^�gxVe~�B4���i��_���2�{
\�ȂO7��π�)��!s�l��|��\9{���\Bb��Ǔ^��$�1rL0#͊���|㇧�u`�lnb*�b�_Xi/��W? �ɟ��դ��Q0(��.��ߌ�Y��+����"�T� �G$�_�����(��?���;�8"�^YY!th@�� ���o�.���;@���w>��ddX�RN�|xb���Ce�����)}"�Z��[���&�wx8���t᾿8�^�u7�Ry^�����Ւ%K�q�F�`b���IL󋵫(ʊ�&$��S?��-z��7,�M�f�K�}�����ja�L]������y}�,��d���_��=�"�����;g�]�`^z��&M��իW�W^�q������}��u�ҋθb���81ԃ�is��.;��[3f�&ḫ��t ٿ��a�_��0T���|����GĢ`���Xw�5q�Z ,/ ���%�(⭷ފ'N��^Y�?h�����3R9�,�٤b����iW#PYw�q!�$�y^D�F<�����N^�������* ��9��}�D�y1I֙wAIg��|��Çg,L̨�z�>� �}�Ylݺ����� �������r��%A�}H-J&�B��6" ���+�2Qpɡ]0�����������$�������ʸ�������^��1W���O��{7y�Ռ�=*V�v��M|��p�u�aӦMhiiAdd/�
莖��?Q1���^w�(v�o����]�U�k@�j�����'pD�y�~.�Tt�����<Y�%��)Y  m�|>�����/�CQ�����X�{�ʕ�o�C���F��;Ώ!L��_��W3Pv|�ҥK�x�bqq^�o2*Ƕ����4DWռky:�p]-@�r"�Փ)T���[�d���ȳ��e�Ć�#�G>"*�Γ��c:����/$���6a۱e���V���P>/�̫l3�׽e0����j�cɘa/3䩧��}��'~��qH������`O!��{ёX����Q�wg�O�0f".�_"�'�B�W�fb_I%��W�z/���Y!�=��L%a�/c�`$"��\����(5}����#����q��A,�U]�s����\/+��'0:::��}c���y�Ν;��ى;�MMM�B-?�c-�;���|3�o��!���9⌋���c=g�m��<��C���'��|A
�|�39�����Sܒ���c%MzxLڗ�!X�Ӯ�L���y�'	+������m��^�X2�P�����Rb�Z�[�l)��}6)(1lmm����E�6}�t��B���3-�j=n����(1*�/Dέ+u8A!�@�<V�0/jƹp&���y.�������=���b���DL����_W�� 4u�Ykl�'08R娴 ��ɁJΡ�l�����K���~�m��~1,	���V��LG����(�9�`��1�uK���aC'��v�?��%�F��܀�X�{��W�O��8|�E�r�N�X���r��*V5�����(����2��xy�D>��+<H�?HS6@�b������F0o)��Zk��7��zWW�w���W��e�������U�V����?Et}(�3^���{�?�)�f4��Ť�h��
��O?�@� �����&F[�Dno�ɞ��QZ�`�J��)J���Əo�����RJ����.��vG�|��$�!Z��CK�)�{�^�Ϗ�	�%�?BZhT���|¡��vv h�"F�<3cjK�T_[�%+c�&tM΄�\r�!z��֭[�K)��B���5E���Du$�
<���ϕ��<)���2R�5���m��Z*���s1ip�0m�項�>zwG(�����F�wM���_�� ( ^QCyz�_�:܏�s�GI���˿s�E!/O�9�J}VGʭ�RAʦ$E�c ��2B���P�$ :)�kD8L�%��;фCgk��hau�@Xt5�H�~�}oL��5R��Q�N9D�����O�	$Y�t��	E�`��E�o��R�]�<���p�]� ^�Z�V�yoϓsb���gw��=vƫ�[@
���6�y��C��&E@ƙ�0Ǽ���b�    IEND�B`�PK   ��X|�K�?  :  /   images/7720185d-ee5e-407b-a613-fa89a316821e.png:��PNG

   IHDR   d   9   ��}   	pHYs  �
  �
܄߉   tEXtSoftware www.inkscape.org��<  �IDATx��\il\�u�ޛ�f�pI����Z�Ց-ٖ�ڲc���I�K\$�Q4��-P (P)P�E�.H
4HlÒ�8v$E�,ʶlY%R�(R�D�����3o�9��g�!9o$[4���{��w�=�|�|��G{~d�KY2�`��)�� �"����P��uݪKƒ�%���̝D`j
��~�u7�I�M�]*�2:;��D�����ї�R��B� *J�v������4N�oCGo�f����.	�ޭ�Kg14>�OT�3^���
)XZ�1�z�U<�3�U�iE����3qT#�V�tb"���,i�D�&.�������E*b�|0��I��	`p���,a]�pg��!����BtC`�m�6`7V����-C�if*�c�bb�\���z!MHhp"�r��H�{��
����� �*��5tNQ0c`�5�^�ċ�P�1(�˚���<-�t��@M׈�;VF�,e,Eq�
^��?��%�y��D�k�aM��i$����JSt�a�2|�q��Pmx���g"״ӿ�[N}��Σ�|k�RL�cMn����4a�]#
&�2�ۥ�R���Il�I�aEg���5�����2^��C���t�{"2�aG.��ae�A��!fϞ��XQ�c�k?�3�}.���g�
�4X&�NI�K�"J���b��t��&�R��;��G�K��v%-�[L��P\�ώ�νF�RV�㟞���������t����`��l&���S��b��!c��)'��<�9H�:����;;�
��'��	���4u"m���������h)OQ-�M��5���^X��*h����Z�[�YL��W9��j�*�P�q�
9jŋ��s�b��l�bN*�P���7N�|�iK'�,^�1�YH�ѻF3c�]1|go[v~k��Bow+j�ޥA�q�ݛ2+I��Ԁ�m�aˎ��E��wI$��#<��KU8N�#]�9�I�jX���vʹ��>�{<fj�2L�<�T�M��dv�h�&H��#A�UB
��۾��i���m�e!`\��cmu�۰������u��`o�E���dn2)ꩨ���_�.� ��mD<Dc�{��U�����=8v��(�g���}^Ϻ�$+������+gttk��ɻ�\��
	M"�c�c��ဒ�����9U&XpzsnR]^���,M{?v|N�PFZ\��T����/?�!1N��D�gRn�E��aB��5'0��"�N�yv34��{���d+ *�
*�3��i�΢���ue؋{z�q����6����7��y����Q���KN`3����ښOBv(�TB�+|��~7�d\�"�o!(2#�))��)!���V�M:B�UJ�	K�-
�П㤐�A5g`�tT��,q@�u첏½ E]����Hn�8r�,ǩ�Se3=�._8�D<J���KU��S�h�&0:m@^D��������*=+
ajj
	� �{4�SGhU�&�I�y�J1S�W'�8lB�h��ب����k���d�v$PS��ehtZ���M������TX���xh@�H�D
�)�G���ĉ>����-��b�ڵ��|���J�m###���C  N!���*z&4L�;���x�xf}?�]+GW�WX�<O��t�_<�]��?���-C(6���BD�d+z����eӕ?�BǗz\�4__�p_�B��HsS��-���|�rlڴ	cccp��ęFQWW'��-f:0E>����m"�Ǉ8�k�o`���	VJ���4�cI+�݄D�mu,�E�ɑ?�(�cm+��Qz0�6\;�{���t�Đ����-�ᩦ�===())���J�Omm-��$�_��r"�_���˧u#Fn�Iq����G��c]d!㷰B��B>�S�ô���+u���"��-�
��;~f��RyL3S�笨��*�"VIȄ˲}Lf��>�-��y,���-��iݺu`ٲe���Fii)z{{��S��W>�ah�1�-4G����:L��2�[˳1�0?�KY!�,�{�yrg�oI3u�1�ߵ��H�ȯ���g
gz�Ǉ��Jh��h���,� EF��Cn��C��P[+#�e�	����x�^7^=��gs���0}��[��h2n�K�� '+�n�O�v�s_F!Iz���d_�w<�zb�}�m�L]�i�N�6�H�{Las�^��� Ɖ��6����k�<(X�a�G[��[��G���J�N�P������V�s��w%�򦞇4��xd�"���a1��N}�2<ͮ0q�0�g�:���uS��o��u+7 4=�}��?H3u*�wm��=�"89�r1�X_:�7^�g��w�OQ֓;��`�|�H~�4MDSl�7o�������8�����ֆ������7���12�+�N�^�"9|�Sز�A���Ng.?���(�k��.�6��dX�]��,n� SO9z�B�Zue��ML��
�Z*k�aG����QgX!l!�HD(�C_�׋���crr��� _f��=A�\��S�jJ�������8�C!Y
�����"|(#���f��1����꼈�k�S�L�cS�<��##=hnj�0��m'qc܃��l��pꜹ�G=@/����[�X0!/��8����Nu�YHj���6b��~�r��5�1�:������
���_i{l'��'����c����'���^���:5��76TkH$����ԯ�8t��^��!S�C^?�6�/�J�I��V�&Z���QL�y��8m�AUd'u݄�2�IHM�9c�sb9�\1���}1���
�Y+���0��j�I���py`Sg���i	)�E&ON4�x(*���[&�$|�a7���/~)���+�[<��':El���Ԭ�v;��/��,`�R��U2q�����~~<���P�c*Z����J-h�YU���c��D	q�x<�Br�z�L�%��ڐ��3�d��������D�NP�rT"��f��g�)+�7�o�:E<$�ȋ�iO�_���}x�)k開9R���W��/�"�W�`[(J��
��y	eqL}v9��CK	��pTGRـ{w,�A┄�R�L�a�(��b�R9��K�	�:�6��J��On(�����GX�@#���rV�
�#N�i{��	P1L1�ojM=�ZS�����L=.c2$�f�	�&Tl��A���B1I�[�DV8I�W]*�NqD�˶�C:]j���F!�n-"i��<^�9_�P��!���{�o��E�4�#�p�e�S��1�ƎSϾ�"��cxv���cYL]��Գ�f���L��HX���������:I8�lI�5�ۚ�輢[V$���"��41,P1l����f���~/3����w>������ԯ�2���'��u/6m���k�ޡN�d�y���b�|F8�L�*��ܚ�+�HQ�dV��n��C�h/�:�HHs�a����k�k2L}3��(9 b�W�0��-�^��.b�!�L�s�8�S�۶4�c�T�d�آVYsNx��2w�|9�n_�L�o��ϑ��\ԁ�ky���p4[T�$�ߖ���`u����~op	Υ���L����i����2�vb���[.���b����=���S��@r@�_CE�,L���
c��7e�}C�K98����:��U�~�>`ny�,}o�v���כ|8�❻�A�v��L}������Ś�ś
��2�O���$I�Sk�t�8h���Z&�ԉ))�F��b%�����u�H-E��l`r�?���@�8��+�x�`΂X���y)�����G�ig.o����b�gM�Zs}�\��X���kK����<�� ���_>�)�����^b�.��6�:��{\ؾ��
Νw���Ҏ0Qt����M~�+6̵�����9#��w�s
���8#���:�S��[T�� /\�A�"��n,%.d�s8�o���^��=��lhY����cSm��0��8��s��FL�� ��E,�k�H�N��hO�����
�Iۻ6D5)��k����pb([eN�����VT#��V	�,�ld���2����sp��㗼�-���n���`.>����d�G��3	9�MvE�[{��1�$�^-��١~����nii��ѩ�HVf���Q����1�ӓB^�3\\)��"8��L�ڶ�Bǲ���&��
�YS������r03���T�����yI�^���C8���ؾm+zk�7�n=�!3�%�
L|g_m��V��"_署�?B��<@L=7��N
#-<'��`�x�dQ���{��j�$|�7���~�%���f�S@�8�ѹ���9�Z[�DK�V�VcR�?�y����~dsO�J`��oaͺ����7��Fp�_IH�);&���cϓغ}?����q�PTVp��`�W�m��ԛ��X�N�!��$��N�ʀ�s׵y�է	��Gb�w����̄�7{?+�0uw�
ce���y���bY�����38�:��L�骚����s�wiy5��F�޻o� �4N� �b�ǋZa�g���c�<r{�����L��X�ײ=���X�ǩ��Ia�l�h:wDN�M��H���oR�
�n��Ŕ+:�t���5��~�!��r�k��@_O�`�-�^�ev����SoaA��X?Z/6����b�|/f���L�$9L����
���� K��u������|A�;/�?�+-�?I�ra�����v���:AVbDFd
E�o�{��8 {���.�z��R|xqQ�9�X������N�q�Y�������ݬ���s*�e�M]�+]N�r�h0c�Wۨ�{�؞r�盜x��4d�W<A�����Z���ɩ�{��EE������4�Cq1��7�xL�9���|�}�W�'/����mI4u[L}z Y�Sg���GW	3u�a_T�Rbq��è_^v[^�dK9r�*Z�F�BBv��SwQ(������a�_>�tSN�1�����0@��TZ��a�t1E�xvb9u�L'jȖ��}t��Р����z�O���d�c��~��_xɉ+n+�o=�sj�۝ضJk �T��^�S�T��Z7�e1���%���2�n�⭋>띚Y��;�j�o�x�rRXH|$U�)l�7�"J� �Й_T0u�2���\Ԯ��"���;(�_�	5���(w�,j	�{�6���k�/�.Y�mw��e�#�Ǩg�-T�^��b���r_��UYb
�R�8�WKڞ    IEND�B`�PK   ��X��@��  ֈ  /   images/a2085874-a866-43e2-ad0b-af370f9f341d.png̺W\SO�5TD� �H��A� �7�E:��((Ho�BCoI�U��N�H3��	Ύ��]��s�[6��33�Y�Z3��kM%*rFrD���R��	]yq�:pGWwwx��l����,~D}n2x+y뺿���������9�9{�X{��{�g�I3�@�A*/���g�,xd��NG'���z�Q�H>��?�`NT��(H���`(�w>v���Eꝭ!���h���3O��(N��k�Wcclq/2� ,)Q�̪��t��'���M���k���x�_�Ҍ��9�#ūW �G͔���b񟼁D���w���W�/V׼���FM|��o������俿��˓_;����wcD�����i����F�x����mR�-C�T[�,G���Fn�7Ū����=1Wð��pm�~����Yj*�-���ҩw�X������{F8h.ӹ�}o���)�q>m�YG��G���5�J���W~�uP�|�_�_~Pf�)���?=M����"P�ی���C&�ѩ�ӽ�M}M׀f+~�ߞF�y>(�<^&V��==����fΈ\��Rd=8�h�2������W�/H��X��g�{;!��h��=��X�H\��QZC�Pӿ��o��i�:]�3	X�|��x��q�	h����#�.��nl��ںY��ۤ�Og)hF$��� �/TJ�v��Gf�����rq�vJ�R�y�I`���3�*�z=5�+Yͯ7�I��L�sD1z�Ё�������� ��k��Co�����M�����ޫņ���8Ϭ�����ps$�_w<&j��4[�J���f�j^�5��]\�`�:jȚ��j�7�}�t��2���JC�ܖuڏ�vEOO����O\�`le#D�5��s:iͩ*֮9+�q�37�d6A�U��cMG50��Ȣ��r+�9r�~?횓i��U�H�G'ŦW:J�~�ˌ3�2� Ο��}j���	~Y���?\͘��V,B-,��u��FI�k;��ޞ?/���hz��F̃�ŉ��!��w%5(�FI��� ����`8�  �j霡)/�Nsi3O
}�!��k�̉d�b�
a1��t7����*"(@��	3����	��6e��}�X���t)��V1cq�e;��I�	�A�<#����\����Ĵ�V5y/r�)�l�/7��+D����cPf�e�g��f�YO��]�5 ��ΠjO��U��7�y[ň�
h\�T&s�]���-��Z,�WR��$w�HA�O)����"���Јԍ�+��"��`��z����U�9;#f3�Ĉ#�&X7��|�%H)�77�#����<NA��\�7���O/��6Ź�L�2�CFBT���;�G�;����4�O����������;[B��N��ݵP.�wJ�r0�z�ݸq������|����3w��@���a�-(>�]������������2/��h�����_���]B��Z/2g����@����ۤ�-����A�	<n��}b
�2���i�؟3)��]3�>�>:�b��Ky���($~�-,�dv�%�ğf���l����GT���@�����;L��@���b��x�mp�[<5Ե�US���H�3�ִҮ#�ڗ�,3����w+�kT,Ѷ�x�Ia�h�=�l���7�Q-nTZr��_ߝ���)�i+Q+���E�v}$�g��\6��1����[d@���c�'�w�3���4��3�K��<Q��C�iD��&kel�;Wh&X���8x��Yi��k*K�����껅�5��\��!���ٔM���y"f�&俩���Q�5b�e3��b����X��/�~?l�	�~Q����{�+���5��'%��E�)�|����Fb$K��>"���}��~�3j��i8����속i?��"�k?���Z#dވ�)�]�`odևX�خO�����L�r��d��1���?��m��q� ��0]����W3�[�����7M��Q�����\�\�w;'4%Wƙ�h�O`=e���Z6/C��ݨ��H����g!���W��� ?���}|���ܼ��BpS�z�4ҸEmF�ٯ{V����7���I�4k,4T*����B;��z�B��Ɩ��D|9j�:�q�������������ҳ�D�&�/6��^��I��m�B�,K�͋igd`x{6-'sj?��u���5�*]�o�YH��,���6Z��Lz<�Ŧ�x���WJ2<nB�,i<���^+�WJK<n<�L)<mǳ2��An�,���q!��o�Б�u�Wk�Ğ�r
����>�01���w�x�?}�E^��A�+�V�m�臹b��LRP�I��<��+�'sؗ�љ/z�0N}�&�4�P�e�(��x΅���Er�Y&Hڡ�6w#��n���a�����zv�K'��˕v����̩�����sE'ה�?>
�9��&�!�O��vL�-#�M�R��+�������zm�\qBH���)o��v]jv-Q�!+V{TΖ�J�z9A.�����E���Edܨ�-\��*��q�M�O�W�F�0���C�Q]̚-���B$��������L`�!.}Y�4M>5�
Zb�Ub������V�>�s.�)Lx	W@��h����Vϰ�&P��z�������Rʷ���U��q�Z��kf��k���F��{�T55W��OL��9m�������H5�η�-]J�.�t�D�@���ݪ�9q�c1G��X�n��t�BO�79 �a0DW�e��+V�#���s|���c[5q/�@n=�ŇؽP���p�P���E�b$�%�1Č�lo�QHN/h'��8t���D<��a�]�dP)H���넆�}���������h��, ��0jaη؜�����ԡ#�҇-R��c����ojFBs�9����R�ֶ��NڤubA�rw~�Py��l�N�	��v�a�{>9���X\՗A�[�@�����}#U\_�+�4�,����7[�"#�Rv
Ȧ����⋭q�.��p�ϑ�Jz��c�Ve?������R&ΰ���I��\��cc�?]�ș+CW�`系W�����������Kf�_i��S�I�K!*\��"y��U�篂(:I��d~�V|��?�>s���'�V�g��<��w�ش��CH����߂I���`���-�Xe���,�'U�F��8�鶵��*`1�d�z�����rg,ǁ��\���d6N��A���Y��<��WA;��-��4�������C��rLӌ~k,0]���{��U BÚ����z��m]#䐐�I1K�$�����k��m�
}�sgɳ��ug�Sn�R�/e�?EQ_=W�.�+NC��_�)���q�lf�F]���Ms���(d�2|B�q�A[��6��(X�����'~RL�Z%��D�h|pg�� Ձ�>�z�x�+��n^BB��0Zᐂ�)�����؜CΫ���X�rK�dA_�R�aa�c~nT#c��dD��P��w5��m�!�T�!;��	iN��
W���陘���4M�W�N�sq�{���f	̊�d� U����Y�_�������~ST3V�]�?�ŔE	i`d�]���և���'ǜ�:�f���;�nqԬ�f�O�r�V��L��A8>*:�0fV9�v�B��8�P�w��wXc�4��N�ڵ��>���ֳ�n��_�������ɨ���i���� ��.:��꒖g�$����(h��~&隕���w�am���^�j�9I(�8�>N��L[�6W����΅2|(����ܦ��Wo��K��LH
6��q�I\�x�X�DM҉�<�'�mk�wmC��-U{�|�.�:���z�E��L����~߿μ+��u�����]�7��xQ���DF�r	�4ҞV�j��!.�P�8������Ӡ/�?���w�PҮ ��ݳ\zC�}C�ܵnË�iMY'�8F5=��OU��� ~�v�FN�3pl�<�����,6%��!�X?���+�D��P�VC֚[�w!�<�L���hTg*v�X�k>��m�2�:ɏ��a��K���ƮT�{C��h�:1QY�=3m�i�o��e�m���'�v�Bb>� )Ҧ��`%�z�N��3���hXO챟1�f���R\��Ԇ���,�g��3��W���j)Z�В��ԑ2hʆEYc�et��VE�j�!k���oIsO�lU��W�j��~��^�t�D}����@GĬ�����������,�}j>�4�w
��>jvNyY8ug20��ڳ*'�=�VC�ưۍL*�Z�F@�<~��3���N)�pRص��G��m1�
�a�M'ud����[{�M���"c�V6MB�ɓ�l�P�L?����?�Gϰ�<!����e$K�	\D"c�h�8?�q~:H�qq��0��I��Tʊ���|�@�+ 獸����@�`u]���:o��"��ݚI��;l����V��	5R0�}�i�}�(M�4��wΖgN��l�An��Jq�6�7�V�^N���j�&�����\�A|p�~i-~RV�Z�m��uMriiQ�u�Xd�d�����ː�$��A�$�����ee��V�W̌;�A{Y1�D�8~y�{�N����c��1����M02S��6LquW�6vbΪ�5e��`7[ �إ��?�*�t�$�j�D������'�Ӆ%Gxc5tz���kN������Ͷ:�xxX�9�Ji�O����c�d��g�UM�ٰ{�ro!,0��n��iB/y$Bj��v�hx�v�wz�(��?ג\^������qf��u��j��l�׎ ���"A�l`��aߐ�󥯠��w7`��%-�V0/�����o롦%-��΄$���#�B ��Ŷ����r������q�S�T;yJ��ͯ������>,��*M�op�T�צ%��CM�&׌+Hw��n2�.��9��~��$�I�Z�ʋi(��Ғ-.[�mj���6n���T��Kb�V���m!���}T��CM%؇�9�||[�������Im�2C��r�H'?�9Ƨ�'՚z���۸%a�rK,�4�_`&���d��~ߏ8^�
�_�"D��������3L|+Na�SL�K
ł��b�U��|�l��A�'G�Jq/j"�0�L��i�	��B-Jo0�Z)�x��έ��S���������Vם�,���ON�>����h��X�.��4&�Lg�a�f	T�0������I��Y�E�t�v��8��v$!����-�ᅲФ���0zyj^eZ�M�"��ss�&�����l�M�٨����y�ޠ�,N�Qi�[�����l�k����e�Ί]�>�]h��J]l���c���ЩZC�����9c��=2aj��}:�4�:�>�z�abی1�"Q
,��<�hbY�E���hq�yI���g�Fr��Q��D�'�Y����IХ��L�k#�~�f��q��#�"g��lAH����c���p��yչ)��Yer��6ηA����Kd�Z��փ�{�[Op�"C�NĐ=�*�>q�����R��DI���頿�M5N�.4_���J��0x_TCx��'b9�P�br^I��s�$Dx�U0���q�}�f�|�P'#4t����v���/g��n�s5 1O�Enz��V���#)���)Ά)r�����`p�}�uҠh��T�����4���+	<����&��!<�t�o<�ĵh��;_V��h+�` ���ΌR�M݉�Z��"��V>�l/,%TW$��:sb����_,�q���֍�?��h�s���H6�;�Z���J/b�3��2Hs`��]��c^~����rI%*��]c�b|`%�
��x`ó��AG�"m�~�KÛ��ŜJ"B2|��U߉V�J��N�9�ݦjxV.�-w�Loڪ��t�]�dֽ�=	h ��+��$��Ճo�"����=,��%��h�s��&j�&��0�%�:T��,]k���R][���}3oW�2��I��&�T�"ؘ1zFd;�yQ �ג�E|�0.�p�ԄN��4�W���*[�a��$ ��9����*�Qݱ=%W�Xz*Ef|8�uIq2�zDU}�����3����p9Z����or��p���=�˯;`�a����<��Ţ*H6�)�Q7S~|[�#)��C�O/�+�g�p.f	�k*[Z�|c.?�&M=m�:
��G���@V��f|)iie߿++**r��"[��f�}�[���m��߆��^aY�J��V������/ �sc_��Q5c��ޮ������k�ױ����A.#��e���0���?�;ay�5m���V0%%eINTF���M{|���-�R"	�C2U�� 9q��_�Z�HV���v�Ԥ�7݁��Ӈ�\�	�Q-ᦨ ���Et56z�F����OM��742�!H��~�:���0�ʛ���gh����X�/�V:K�]vD�w?|�0iY���1�ws�B�L���c	�1v��b�%!�'��T9gN�!tֺeH�HL���uSr�[�L��	؃���݈<�=N�J ���"Evvvch^u�k)����
���ɂL1����ؠӭ�QWRGC��or랄Ӓl+�p��x
݊�\�m�ٵ_/�toz7R<�Hx!o�Ԃ���-,�7���ᩓ� �=(�d�|ǟ�oaQKM{�n! Snk�3�,.fu�����ew�(Z�����Q�)�pX��Fc���t
����T��kنC�R�#�����wد�;3�-Ԥ�3J��8F���'��)!�.����9�y���Z�d�X�<ǒd��黽�7JFZF�'�~]�}��?x���;�@O��O��bYJ�P��m�����������Q��š��������jj�::Ӝ���++5EDD0[[��x���&���R2j3-Ɇ#ߘds��v����?�}�.7��Sm(�������I�C,V�d��릕�K*�t�;Q����ip��9���ϕF*P5D���u������S��@&�W��ny��UFVV�1���3}�⮮h��6vp�s@X����3d����������$#����&�dpppjn�a=�/�;/"�����&f�����xxL
�ֿv�Kρe���SOP�7��<Q�Ȍ_�k�*���P�Ʃ*
{X|��I�vS�d�!i�ycde�n	>��wt�zd)��Y�)�ZU�����䊗�BxTt�nS�S�ɹ�oׯ_�B"ˌ���=���X;���f bpt�ңrhc��Է��:B��hN��+��L��FD߭���������^��RȾFi�@ޠ��6 ���i\i��,�}���""���<��{&y@&�B{u�2b���}�f��\�$Xt&�#/u��0��Y���Jy;�M��5==��
>yt¿��?s�~������mS�K¨�+_r��ή����֤���^R��\ԫ`§�3��uu�pQ��NR�k��Yd��������U"b���c�?Z`nl����m$��ȇΩ��cR�^�W�>zu ش`��a	��{�;sy����!歁�II��U9ii%}l�f��馊g˃@� #7�-5Ӿ�l��b���n)}u5� }��=�̀@F��ΆA\L�ϳ /ٖXgj�B4��w�H�A�5��zw�����S��֖c�ߕH"LkcR�[PB�		�>u[�sU͖�����;��W�"��~7��ݖ[���H�{a����Ey��xS���1�F�Z195�n���~+�	��[T�Q3��J��cSx�ޭ�>�7svr�ɖJ[b܅TV���n����s����w��j��;�g�1�!2�ul :{�[;gX�-�����)g9%�n<�y��*qR$�xg�#�����"�aճX�j��N2��=�651Q������+� >�m�_9�]��jDD���ܳ��:��[$������%&�GU}���	<5Z<<�$���b� �_׿~���K�nF0�*��#0�2�)�舣�=�lIU�H���ӡ������Jss����S�)��6L���?X뛞�o���X�iB���WjO=����|?O��t���S�����\y`\fc���@����/?�{�𹩩�{�7���6���=##� (�[���������h\��[t�
�b�8i���(腁Jk������s����E^r%��B��O�7
�gn���������LDm��QO&ho\;^O��c�����[-�Y�����YFՌ����D5UU�kǍ�ShV����\`���"Z�%�i|��o� �@���fD�)��\�Y$�Bm�/̵ָ����PYb�Rwɹ��]�j��޴���9oprrJe�A��cW�]���g8'2QF������4 ��2����x�3j�`���3��E���� 4�.�9fd��k[[�Dm߼.Hi�<��Fa:�.�u���h]7�''v?+zP��"��7���JfX��%����;�lnV���|��o��ӱ�l�EH3S�LEt�	�\V���n%�Kz��3�O�FJ����^Td�y0>�PoQ}G���]zZZGo�㋚�8S)�Z���Q3����R=cc��ꛀV�8������T'Ұ�1��W�R�#�R�!��VM���4]����$��S{�G�kS�W��ͤ��N���:%�"�
�������a�t߼�����,n�9�N^�g�ԛ_�H@s3pW$]vI�ޢ�7�'��Y�nv�O��/��k=����.�ږ����ڨA3��)��ת=�s�v܆�V��0�
�=d6/�����395���-�� a��p�� ��9t����|q�Ν��
�8������|��Q���r-�_�uw��Ǧu�w�kؙ\��̨V�Fn%{E�4O��&���p6����9��M��J!�`�;��L�Դy���X��n�ͽ_�W�4�p/2<[�3-
yv����|7H�"p�������Y'#�|Sçk�9Ms����>���[ZT��{��� ������x�(�qi�k�/Oҳ��J]�Ѭ�:NP���|�c�d�oW͐v�"c���WT��}:��������6S#_%y2�����Lz�̌�	 ��s23'���^����~��Ξ�r����9@�ۦO���ő������U�V���|p;�je}�H�>C'�Q�N$��m1Wk�p	�򬾈�t	�̕;Z)�����ǓDT�ػ��bOb+Z����/7Y�|��TZU��P\hm�ņ�M:;��$��2����ͺ����ֹ��'nS�`Pz�Y�s�o�l�^.���J��d0��Ч���ٻ�3w���ڦ��PWw�����V,�6o�xN�o�Ҷ������>��77�jco�U|kuV��c����K�~5Ӑ���i[p���m�xZ,�5��D���?�{��vo#�z�5�=��rOLL���A�.�;:�~���+���M�$�QCs��������#�ۏ<����l��jlm9ﺕ�Zxс���zC�N�)��֙$v H�	��5O_������v�R�9��T搖��q�Ѡ)����&@a�$�G|X�Ŧ&,(�ld��S�����e6hr��MM�C"���gs�� T�����!��Q�@�'�����p�}0�y
���)�T��n�B����� ���pM f�H+NN�BBB�P���v�'����V�����G�("���h!kr�8�]���\hFэ$���������=t��S��>a�з�ml��0Sػ=[�/w�,NF2���K_$�t麅�݁OZ�(��{�"���sNx����SS�@���|��n%޿D
|������q�� �.�^��WA��|ek�*���-w��h�oqE�a|���Dwgg� ,�VPb�SA[[{�h����n�+]I��96b�̞�ܣ�e�M"g�F�3))�g��Q,����[G�o�W�w��%����m]7g����/����S�PH=�
�k�r�L����̅�e�	��IP�����!�	<ʾ�#Yxm�yG�� �p�=D�1t��HM��>ۑJ�YSo�o����I+{� ��f��̻����Yʪ��P�[{Ҹ���3�����nN������ଦ"�_��S�
�a$`��)[� ��d��h�A@&L��K����H��0���� 6Sa�h`ut��Gf1\VH���Ѝ�(��I��N26@n�/��P6T	�h �-�k�L4�n��y1ӌO<h�����P��w�yuuu�V_\\L��& �k��6�����#��4��~ ]�ЙK�*��A��o9�~����Ф�M;Rj����͜��T!�+�[���g��� g���&1o,f�����^D�̌�������J����o��-T��2���>FF���S����RDp?�5"��C���;�d��:Scqo���
d���KT�X�@!���L	���w�/�Pg�^[t�7ng>���Ą΅qЊ�2F�o�wI@a�5�4u�f�ַ~��������	�Ɖ����f�0���X��^J*M���]���^��~���a}z
��)�K�o��?�x�yب~*S������n,C�qa����B]��&6F*EX�|#� �K�LYB^�%jB���}�����3@�24�-.f�M�������:�/��R����`�3B`�%6|��V���}���`@X6�/]?^��3>r���V��o {����:~w���]e��W�5Ǟd�����S���R\�7���{34��͙<�U���Z3n�Gگ�Y��YC����3��	њO,�����[	|���
�ݻO����O����w�*"2���Y�4+�@�H�I�� ��JCU�t�cgM?��64'���d$��t�*;��q[�.��H4���,1��&�Ў�k�Ɖ���p�Z�`d#�K�V��m�X|@5*��2Y��("����y���3�7l�2wW�1������405�Ϭeq���Oލ��5�V�`d����	��nV�Ջ��F��\��ųn�u����uo�}6�ǷWK��r�� ��)
���rX����u[�T�74,Y4�f���1W��e���`�����g��)�6�����fԕ�,n1�_�?��y��\o?��S#"��^���{��B^���N��xI �fe���s۾~�h1'[�]����Pw����Г#�-�(a3?�aD<��X=hP�̚���Ȣ��颍-:W<�~(�/���|V|	�Y X�"�e��9������F��^?�th�Y����f��߾��x���ԡƃ@���[an���a/��e����wl	��c���ɒ�j�.gr|"~g�Nr�y��I�^A�"���(�OR��=�["h=�_Z�}��\eX
�2�� �H��V�,v� n��(D� >كy��
6n� ���+���6�2F,'GG���hkp>�yv�훶Z�o�{��^F��x|z�r��R��1��W�����+�Y	*|~bő��g�?u��zO��.��I�T�&{�@2x�MZ�%�T����j���~GP���j�>>>\�ԣR��O.�SMv�AѨ�����B�pJ{2���C	���v�1��|���Vnyxv�����	V-Ҿ�`Ƃ�.̠���25;z�{h���zu�®�� ĥ�o�Q3�vt��LDD�(=��Ӌ=k��o��Y;8k=8�8
l5���;<:J3W�c��47C�[ZVU�"L�F�5��C�; �K�U|xkHᜤ�4'D��8����+M��69�
��{�c��vp���s��b�^�]X9L��2��D�L�ō��B�;��]�)�a��x���:@�i�<x�̘��)$]brNNN���F�'
�� }�V�γ!��w
 �P���5����۠0Z�n�a�B����-��CC�]�ݧ2�*��8M'wꩌ�>L�]��4�V_ŕ�=/$?�U��9�}��w���Q�/�%`wJ4�M���%;$�[�0"N�G�;�<:"Q
 #W2�.�����7^��jm���2�zگ�L���bN�X�>���ëCv�]���$b��pI�Ü�W}=~e�q.ퟌn[#�=�ˉ��,���/y��-��?
=kG�{y u���d�EW�`�0I����d�v(N58[��]�M�on�3�*��D��3��zk@��|�o$I�N�~ky�s�v~�i�!�S���F=N���Z��	���Sup�N��N���q"]Ȟ�<kyb"��Q�(�~ww�.������^*�,,� �rʬkiM�|f1z���R�v���E�>�w�߄��V��քߴ"6:��K0�{ZZ���x��'ѹ!F���&���v*ï������?�,k�Ov�w�n���a����=�ezPϒ��t��2��f�lS��Ohkk��׷pj+^�u����s��g˗H�`�B��d�P���ڻ{�+����	=��*�l��x���xأI�{�B/ٌ��^������%�w��}��rثg�Y���ۛ���^*�����"����F�,bf�@V�|~�$ku8Egd���R�S��\�[i>���-���F�U�?��)B"� ���g�-^+���������訨u�2K q_`�H��3��z��|�{H���c�%����å�%������ξP�8��~���a�C^�s��E��.�j� �7l��Z��"i�*�s.�C>7��h�m������5�)���ه����p�В�$��� \�39�>�m������t�Y?���b�!ٕCp�j�ʧ߿�%$*���pTQ�؞��P�����ga�G�b�
)))��=q���σCC���@�(�c�h���-,*c�T�SZ�	�����)�e��Y⻿L�؍6��k�}�Y�W ���>,�񨚼�&�qnշYW=�[��g�)��4ۿ֚���j�����}��e��Y�i5��`�[�M����g�WG���>�ճ�]���
椄�'�����
�_��~Vh).^�:}���#��֯�������oa�L����Ɩ�ؼ��u�
�?�g��l�<::��lLOM���;�qjf�nedbB�A���b�,U�
�/|���ʑ��f#>3�xJ�m󽠜]�#�QB�%�
��J-����z���Й�f:Aʻ l��NhZ-ط/��Ϝ.��{(q�z0����S�[h�U�H�5W�ǎ+��T��h����%>;�G��?��/�&+K�����~n���(\�m�� M�^�%&����7/ ݎ���wu�-5�:88��e�=T{~D<��b���9�j�ʵ�8��� ��ڣ�%05�gŖ�m�{�v��gg�LI�1]����������G������싴��<��Ћ������'��?^��m�R=L�))���w?�Gv5��&/D%�	�?��;��둞��2~i���J� td�^��N �/�:'��X�uתu{oB<q�BU�G!)��e���d`0`��x暐pp���q�@iu](�`0�pMӯ��>�)�4�M��������p� ̚}~�u4��
��od`K��1�L��۝�������ǈ���+aw�R��z��΁�վ>[>�����{�z̖!}���9��ᴍR{G6N���E�e�A�\N�-D�p�Ѓ�z���M��[�r���:F66�w�6�� � �h���WHN�d�!���d�0�F;{/
j���_�
�������Ҭ��u�,�`ȴ����;RQ�1�&����N�����v�O��E:��5Pޯ)3��!@"2�������LNYM��)���ޯٴ��j���S)����X k+�7�[��9(I�8��H�6���QA}p�R��eG
�Z�i�%�G�81��:���c��[�n�P8��pi_J8#��h�>J��Y�k
w�dy������e���p`"'�׊����!�du`H[�%l��.�qq�G���Ӯ�:��e~��Šs�D�7ٖd�fB��ˌ�.���}��;��-w$A�̌�lsm̶_�$��{�r�]���@(~���?�gX��.!�7�\�)�>�Z6n���;�?�v�*�E�������#���_��x��U�ܒ~�3vxx�g`PE�o`���ɾ	,�X��$|r+�k�-�.��`�'�i�yW�˭�%M]-a�r1+�u�K��S�cD�.g���5C��Sح?�t٦�b���g˽&gp��]|P�y��������K����N6�^F��ܹF]�0숰�RK����NC�OJ���Ԃ���V͖ML����Z�:p�Hc���"�h�բ
H*��R
����G��vڿYSC�Yˢ(HYk���>���� I��B��j�ڑ�{%�ɫ5_	��C��%��k!�q�̤N�If2�)�G���s��Y�Z�+�q��F�:nZK��z��+�4ǝ���a"��U���ů���xX�<�������]f���P�	�
ُ,�0]�oG��Z�&
��7l.b���n��
?���UC��7^B�	R���?q�]���m�(��Z�@��<���짽�F�f�,hu��C�ķ�E���Vt���?��g��.#�`������J]Ϗ�����jèm�&�M�� �w�3_`���j)I)**����l��W�tu����0?��z8 1;��E4t����m� q&�.@��\X���9:���;dD�J�5�c#�VdT�bƒ���[��F���ݩ+U=�Q�Y�D���{,II�g`�~܂A-T���|���]�y�Ƶ��3��P[�:�CVB�@��<,��+J ��E�U���M�d�g8JzL`�њ�e����K����E�f[�sBa�+Y.���=X��hU]0�|���i�>�S?�i���U��:5�B�y��Ex��0U��C����Oxt��CTD��n��͟t�k�s������}I����Q��<^S���
ޢȟM�X'�O��"�M�Jra���{�l���Z�J^�v��$���*��V�y��鎞�>WNv���~Q4R	��q����|��2tTc����3O�{b~�T0T�6�6�b��d�*:��d��@��`|3��N�����h���xlj�[R��][E�Y'�A�~U�c'1���֤�ƫ�r�{��SO�#ˣ���>ǘ���ͱ�Q��u4����L�vQd;�=���:;&��������3��Ĳ�Х�4�����4���@&o~�PW�8�u��!�D�BKZ��n���N�23�5{�$�u��D�$zڋSV[���k)���	��#��B :�/Y���֐��6�WJJ>��1qq��MM�����n~N4���ˡ�����E� ��q�'w�	3�8xL@	���ܟ=��e(P���#5t�aK�����?J��γ�$���*Ô�G��t&g�	8Ε�;_�B��jl[�a�����Ҭ�P�������dzZZ������,��(D�n��Ĥ��1�1-&(�O�^�X�hj��@ܼ�N�w�;@[eA���o�)�(Ұ�%I	-�0�W���%0)�0	j}Ǐ��u����������w��=�L�C���:9��ܣ�&WWףX,Ƿ�?*<),".�����v����(@	�ȭy��m����ծ�@���
�	*�Oe:|7?Mh3�����-���D�k�e���0��� 	}L� �҆0�1��-UW~+PYAI��3�� r�Ц&� 7_�g6 �ه_���l �HlSss���?YDMKOo�D�H�d���f�ʯ{� ����f$R$J���>�=��mA��f��,��]0L�閞�B���x�O�wSS�G�w�L{\�H0S����&�����-	��C4���	����w�{�,�������3���w �E~��O�i+..~� �<�R�6��Ի��g!#I)�U=�§�8��d��(~���M�l���(���΁��٦t)��d���<��J++g �Й�.	kd��{�컫���08���#+�LGG��6��2���a0}�18���Ζ�ُr�ա���m�c'�Κ�Қ�E�j�I��6��j}��ݏ���:���!W�v�_!r+�b�d�VYm�aBw{�@���_W�;l�T���|v�(���.��{ tW�/%Ԏ�"r[[�u$�ȼk���-SJ�Kw��$f(�ٽL�� �֠�|���7ܮ�羊i��ѻ�=wfCV�8D�PN
�q���ŷ��~��^\\ж�4�lo���&122ޥ�ξD��
�,��S�0a�u��# =YZV�V�G<2�=���٩ר
�uxQ�ydU�D�+,~w����!�/F���z���0�UøQJuu'<9�/Bq{R��gmG����j���/Ku{|�+����e������\
�eq6��q̻�~����2TC;Tkk<����������+W?Ͽ�_<;�H�չ����*��>2.!��~��-�'�p�\\:fI���><m!��'qj@�<Z�p�&>�EJA'.{���-Y�[�	ml��d���&� �4rh��������)�m�WtVa#����P	�;�KO�·5�����
�)W�ɩ��#a��s�P�kY]�nEEfs3ޮ�)��yV	I�}�~8;g٦&��/_.�0�J�Ql��	'�+�0t����$����c�śE���:����
;|ph��6�[��FJII������A�ǎ"�(33�$���5�MVB�I�=�5�w���H.��H�ݣs#|��6W���T�$�k(p%�Q(^#�}B���p+��]!xo�{��1$<E���e��R������ �2�uo�}�7��w�"m�9O6�X����kp���M��#�14��ea�S;>f����p�?�ݳ>3{{siB=.�F����i�ꚸQ��"ȣ�HW��{U���{HGP�(R�!�B%@@�މ�Ф%@B�Kx����Ϸn��]������3�g�7{f��W�m�N�G�^�>��0�2C����,		�A������~t�^�
�I%'��a�E���e�>ڿ��� Ej�������̀f��y��d��-�<;����Xe��R��z�M�LyE���YAB`����'$$�#�חu�o6y�V�txL��뛲^�߲��W$�<������կ ��h�-?��x��4_x� ��*��wN�d{��Իǀ[fyhV��eu{��8L����l����z�Y�����I����l�g��cSOU��*Ʋ0�-G�Yd"�ϒnm�Y�j� R���Ҷ��3�b�s �Zƍ�-Ve
�?£M���۷I~rE���j(�#w�3�2cA L������#C	?��t���w�ja���snj2�K�K���F��ӛ-Ɖ�%z�>�뜊^�|$'����$�hy�hc�p����+��C��oFQ���t�)��u�}�ǉm��OY��}O���"�* ��z�eI��|����ȳȚs��A�-�?�e��G��X9:�ʨh�!��Z�V�tbς�F�#��
�}�ft�׽�l��㢝�R���D���g����V����b/Ox �i@Z,R���
�8�^$��e0��VG��۫�Τ�5�ȡq�?Ϸ���� �&����5��u��E��	�'R3���'C�b9v��ēn�+Ǭ8͈/K��,��Sr�و�A�Y��6ķ�Ɔ���e�OJ�
_�J�S��S(���[Vx�꽞�G�!�p�;�v����Qtmm��Oٕt�+������!X ��þ�k)���/��5�?I�&�7�U���	0�3W��w�>��^��d0>�'�t=�3����m�����R�n���=n	�Z�׮�_	�7cq��H�4�5^��A��V�7w%�->���E	<|Ϟ@���|�|	����sm���[����{��&p�]x�sk�L���Ɨ�#�s,�I#k�D��m�����ֳ�_���l"E��討���u.*��? Z���I!����U�0��2Y�y��`�>@�3Ic�*��AO'J�d���}J\+��BE �Ҿ��E)��j8t��;��ƈ;6Wq�,�<>��J��|f|[1�����'ol3��׵�g���D���[��CD<�ޟEſ=a�UDY���Ŀ��݁h����ٸ���vZ�ś&}m�=����e�0W�6r��R�����[�|��B6�9����ƛ��K�[��G�5��_����)e9�g10�D��[�D�P����Z���j�Ъ�j�5���+�)��\|:�P0�}��lH�� U��bk��%&��'��)qޣ:�G����Y�HO�'��O퍌�I6`�S���i����'�ݬe��������`2P?��A�<�>1���%��Lw�r���qD�\�a��bA�y�y�'�������o�r��I��qjU � ī>��#�(Eo1��d�C���*_|��6;�z�<���`�ˮg��U(M��{Ǻ@I���S�}����Բ"놨���݉	C�{7x��i�O�AC�3����|1	�H5'�y��Lf����>�ax�ue��D���p�h���)��o�߰��5�ZZ��9)����(b���4�� ��_�j��'C/y���{j4��o[���+F��G��U�A�&�h�ݠ~k�g9͝��~!/kr�o��#�It��\㟺���D��Ԣ��"���d�R�(�w�&�0��C7vǙ� T���'��]0\�}b����Z4MA�G�k@���[��(��ыQ���*L��$�$c�f�9�d�}jt�ć#T[w�ؕ�rDc�K�e,Bx��f�A�P���mJ��G!�����-~�l�\���'�}[#������[�!Iov�@ēl���Uq�g���^$!h3o��7'Nh��;�1e��	�jC�6����n�h;��T�0�%�h7�/ ������/"a���♏[�T��
|W^��Y�j0I�]�T�9�0���(<'Rc&���5�<?t�Ab/̆<Pô�֯K0e_��V�������k����A���q��>nƤc�\����T�:֕#%�Ԙm�s�����G���]2I��� �R�t)�Q0���bk@�0��;s<��/�E� I�,�*��'%۫]�'�hhn)(ĕ��w��^��������L'�#g��fF����^������ظ���o,do1�����(h���M��3�s��oB��M���zƽ�w�T]���K��ܫ�SwF
���E
�ŊQ�FR�K�6K�Mzr+_8R�{[�$X>��%�]�c���<6
��۠��|�l�HbL��d��Jۖ	.b�IH^l��kj��q�G4��3%���)���"kV�,�gIr�.����>XF�愹�({���c�Х�W�[]�5�C��Z����I���_~_XWx�R���:W��2p)��������x����^�k��Z�1*\����I5d(g}������:N~�<�/4��Q�3�+'�P'��	(�/�.����G;=g;3�FԎE�i���a!qUaR���
Y3|�͜X��^�>I���8jq��BCᆔ�ZX��	��(k�k�a�g�<���fW��%ÏTR�77?�+v�	4O���GЃAY�y�����w�Z����O����[��#��Fj�sB�w'����]dTh,��4�x���������#�	9hn��7�?�����	� ���"ړ>#W�l�}15��ͯ����6�mQ]����&�:Ȉf�N�Io� P�[��Fa�ѡ�;�.�)u�@��U���=��6хt� X�Y}��Ȥ�HE]D�Q��"�¤'o�#h�&���V~�������[Wƥ��t�8&�&��U-���u52{V�Y0�7L�Wt~%���^C~#�?��Ʉ��DIp���W4zm��=���4��:�	�(�E�~R�ৣ��B��p4��i{8�%�*R3欳�=���>�Fl|�t�*Y,U���Q���4�)�>嵏�D������	KD��f�r� �]��_�Y��SsRS�1j����8<Ύ���z�7Kה<��:�����'\{�w�j�X]����பb�$����z�3L�@	����6w<��o"`u�TyM��1q�!g>?�f�[�;��������X�Q��m@6ih\.D��E���� �_j�`���3�x�����x-���^�;���������)�������O'y�Nt�Bܱ)vk�8X[�Deo�����{QxW$��Q6S���t\���`���+~ת��ᄬ&�����p�^�I��Ǚ�k��o\Db�8
.T1C�܂�t�N���rF��($^�a˵'i��b��=2�cc(R���;�Ɩ��>�?U��z�G�&�+OJ�ZT�M��Ϥ�Ѫ�G���W�oU���G�N(�{�vHy�b
 ��ڜ����Ь{M�;�W��'bV�[����U�Hb�$Fd��h����6�Y����;��ibF��E�p��B��Kv��)ׁ<���$���B��ŧQ..C����O���w���z�V��d�+J]	�Ǘ�b��(�\಻��4Wq��WUHGǸK!���g~zLژ��K��ݘ��`f~bD�jĶo}�x�S�~��}���z���#�'�����hF���믭Ѝ"�E<�#� /���<x�4�A?�u��m�6*eQ�k)��쓌�6n�f��"W�Cé�Z�`��sI���jHd�DFB%w�����'���5�ޏ�h�r�W���hjϱ�N*@�&k4G�L\��aL-��||��BE4.�,�#�$�;�����a*��X�kT K��2O3y,Vc��z�`�L�`l�[��8?H^�
�ܩ<�h(���"{B&H5S�ϡ��ڳ>��=o4[N/��s���L�3�� �D_^�]='�\
q҃�О8�kuN��Vx�eL�jE��&n�D�;�����ٶ�=X4z1��>��m���G��=��뗑�=�,Qa������������:���<&F��%B�Z/Z�(����/�\0��ss_�=î`�z�����fIJ��+�&�'��e�X�i.*�'ܐ���+�8�>�}"Lv���ޕQ������M��������?�ݩ`k��]_r��*~�����HIB���==�v�\�U�Ӛ�/���C/�+�������م!���yN��Q��3�ȿ��a����/o�ȺnI��A�]<�
�b���,�oT{��f�o������d����4�w�?
�5��H&��"(A?��=�`
������|{�jc�=��-5����s�7%)I*���Υ�d���ڻ�N�ͨ-�'� J�(M��W)��E���|�!|�#�k�%�_�=֐v��mn����S�׹x���(����w˜�i �rS�L���Ј|�N��Mq
�[��~�.�@V�j�#�Z�Uzm���)����o���������I�s3������W�����M�&�2<2�Y[���{�-^G��E�*%W������A/|�Q�|/B���F���,M�C��DH��Wn����'O�l0�-����cm����� "�%��}����h����ml���t�9��:C���a�f;�|K�������峳r��O�L�|�ud�i�&]�'V���c���Q��ƾ�ic��ʼw̛o �&L��)�Xt�,����4�B���ӶY��k����%/ VѤ�M��h�Izv�-�1�9���D`��)��)�L��I,J�4 ���η��X-i �>��T���昌4�N�`��� N��#-e�Ŭ�}�p?�Ap�f��W}��A�O�"�Y9K�>��5��>=�����c/�Q}?;�~k�z�9�nf7(�,�8�tv�C�P��`�5%1�RD�?uؗ�O��g��G��z�r�D���5T�)��6�#�b]�V	�m�4�fgk��?�~@lF�c&�i)U�A�#u �js74'V�����-���j}Z�$8��Rkd868�jI��a�zh��&�_*'l�B	�����a��c��l��8��Hu�|ս�S��?Gި�v��fJ��x�=��\�a٠UMy��0����8J�m�4�u�����az���dKhHž5!�d���V�e����t�����H�Ђ�Rw�wc�`a��A��(\oc���"���{���Y��X����F��n�2��!M��Y��K�Ǎ�N�5�0O2"��
ߖ)�������׊a���X@�pviBy+|a��%�o	�|����g�R%�mn�����)�x�U�V�'���A'0�|#V�;hN�-t��	&
5����-7xM� ���\�`�`0�A��%���u�sP^JBW�*��w����&�`0.���vz�$%Mz�o~�}З.�'wc����y%ó�4(�
����6h�9C�>�Q�0�����d�s�����y��!K�
�c�D��y�a!����kZ����O*Xᘟ'!�P��]����vPsнqeO����_B�Du�)���a~&iÑ�o�p궕���=�r���K�5,,p�g.l���w�[|��Ò���HF<!�т��?6ϰ��T��i��~�w,������Ɯ;�_�a�'��B(�ƺ䐦볖��m�\n8��o#eu�I�@�ι��ҵ�T ��v_(%���)�:��ٚu��G#8���y�}�D%��ƚ���ޚ���5=cY��&�of���'Ak�g\�u|xk��KM�ŋ�7�ۯ�C�������x�Q&�lA����n)�UQʷ�F�ˬ=2m��Y���e��1�E��S����u*�f��n�=�a�cK�V�N"6F���g#&�Y.��/�K�=�m�۾|F���Y,I�6�Gy����,�1��,bZ��A�d�dOV�m�RawΊe��_s�t�gL��V��>�A\_G��^abd��נ3��mG��ޯ�73�웥�(}�Jڝ�t8��.���!#���nG��W��esf��߻r@��*���E����s�j�����h����^�[L����P��,7g�D�4%=�w�{�����&b�{"X+ ���(K!GCP<���eRۅlM�"ϒ��l,�>��T�[,��?^H�r����\�/�����E)�o�z���x�ν�*��:@�湦�˽~��׿ 
2E�36�n�,0ȂӞ�sc���B&[�gI��SN����P`�GVc��]��S��i���>��Vbh�����z� ���@��M/�6��y'�8޾{/��fk�A͍��g&�V����=�n�Ȏ�q������7~�����ҹq��N������G�
�a�f&�Ĺ)�d�da??l�u-.u���� �����3-2��F�}�Cm� A��.��P\��3�Z/s�8?m��o�ZHgwq��l_<���-������/���SA6�;����+��sl댏��4|�=5`�5�|b�����*S�_��KH�"\%�bX>��F7z�0Uf��?aCl�mIeN�d�����!����3�e����O��ۧ��+���VΕ�ۄ/���8D��6� xK��i�T���H��,53ʈD�<�n�&���Y{��)�|��s%H��!�rdyEr����`�ξ��h�~J�H7N�7�x�K�Drd�aR<2	��a�����u����bw=?`�V�e���k�-}����JӋ��f�����[�9���L�<�΁�������+��v�U�b@��� ���`�ca���=�2/�0!U9��hn�q��+8�0��Z�Ø��k�d(���p��V��M���u-�͵��2~�g�>q�l����_g���y�Дұ%6�W}+����5��i����_܄�gc8նd��\.�@��y�3'�1O����ONa4g�哦���t-�X�I�n��+��!	���-�#�晋�$޴��P�����`��L�����XG�'�DEz8��śE��j���!뵀A]o]Q�?�s����<���+ϖ�i���PFm������eb.e��Fn�A���sm\ޥ���x�9pw�a�G�kG�LVp��2�����I栉���R!M]J��_+n�Au�� )RG�L󓂑K�*�n��9�l�'KUg#���GXH��ft%���U(G������ڗ��w�ql��D�udx��׻�e-+]p�2�R���Z,�7�j]}7�]�i|D��+�A��ZH��)X�R �e�R2����إ���G�u��ӑt���T'���Aa}n���	5�4�UZ�Q⬎u��m��RO�{wc?����ب(x���f��l+��/-��z8�02��I]�]��{+Ti�8�W�	6�<5�У����R���"T�Ү����L��a�P�^z����(�Ѫ���|�{W�;�i�S �\��_���F� �&e�aڟ��fA,0�焎$��r�5���$��"d����U&TG}��������l&��HG[�_W�7�I�|�"�6�&oc�������͏Ń(ƥ�ä}�_�n�����yF3%w?A�q���+y�>�m_г�D���UW?��V�V�V�����j^]��w$O����IO��7Ä�Ǐ�3�ZZ#o�r#�tZ�@�e M�M6:��!�Q��J
�K^���݄���J ve|�3]�
�_=R������1���$Q��c;���~mLԑ�s1��chx�>ieӵ��>�W^P��G����:����xpTq�a�[~�����>z��sc":�*�8~���fQ,�Q��ه�D�?��/�U�u�DiJ(^.�+�ikY
�j��Үr�_�ǲ�\e����f=�D��ѯ)�Mb��Í�쫀�k��K�+[-cw�u�J2��#<÷.�7L��'�8,_������z��I���s4L�	ڈ_�YQ����}��2R�iM�J�[����c�I��=q�v�r<^9P��5jsѩX�������AݚK�!(�)��i����A�g�;|�����4__��|�]C��v>O��'�>V�S�wS����,��&���N��?(§�>F*�&��lD���Վ�ܕ��7�G���lO�K
I��w.���$�PO
��y¾�G�r.6�9�9���W��%�*�}�.1�
��ݴ��#�8�P�4�:�,�(�r����̓�t�LU�2H�?t+�mNN�0Q��
�BP�R��M����'_P�l}��4��e֙��O�4W]����"�ErǾ/���n �Jx�U�:=!O%��˂.~GD��۰m�D�{�&G�J%�:LSQ|խ���H�o��r��ݳ7=YgT����=�o�SV�Y�U+��A_��I�@XĢ2��J@�����r	�2�Epײɟ�(����g�m��S�%#�Ǫ�Z����
<�vO�y��;�&�(a����c�{S�h��,/%\�w�T�Y�r%�i�_l6����D���#�4(8��h�t��I3�mzd�D+�$~���әW�W�4`��_�T.Q"�T��b�� ��N�x�\i>�Y�-�P�{\�U�닉ŧ�����_��=6�>��n,z3'���W::)T��U&N���zCoҭ,>��+;����ėx[��fd�c�O$�C�DarSy3��g���t�+-�}9V!8�y�h�i�'x�8�&	#�{�hD�����P��xsoh\��/��#�]��=�%��W]���"���I�3=�Ap��i��>�_<�_�"M�J���S[���P���985���b�r���/ȷ{~__�<|�����i���͙L��'<��A���,O=8�Y�����#WA��	֡��
q �+�}�W�]8F�����`�`���pJ�:$�!4��Y�F��#��'�F)��<Q u�����^�M �M��ր�(�s�t#����z����*L�����о��h�#���"k)�77d}=d���P�T�8�0����b��P��oO���� !��9��%�W'=�s���0��s3�%�芔�O��a+��*��ט�Wv����3��玡1��Uk�n!���H^~�"6`y7���1��AҦ���3B!���2s'6�gҠzmu�gt&�K����6��`Ps@:ݷ��M�2I�r�mԚ�L�-X�P���?�zo=u���2�=��%͢ga�k��+����S��)(A��O�.�^)��E�@�2ψ���DmX �� ����ɚ��LZr���C�G�[B�;��	7�)]7�/<n��	@�����3�(�;c%�4͓k#��^���#{O�WŚRH�R�^�s�=8����g8��\d�$m��o�M��Y��dR�Ϲuv�ʾ��5��Mp��Kx��AR��k�*V�uAs�Ci��_�+F�i�N���Y*<G:�'�����
7S��>�p�5�Iޗ��D3G�TҎ���T���	l�V��������?E��Ф�&��z�|�8vNe�ۭ�X `Q�z�<Rj<���=�	"q9��9Zo��2� �E^���>T���۔�h_��=�g��\'C�  Q�hM����?罋� 	o̇RkYf���Ŋ-����A4��Y��d���&��f=���&����Qũ�,cQ�iaJmE�O�\&�ǣ3�f/�^+7�O[|���5=wg�~��<�w���qF��Ҕ���!�%�k����r�m��4�����@15�� ��Z<�Aҏ��иo���W���yXD�'.���(�=���/��-rwrh�xr�1C��Ay&�}z�Y�jV�>�8�ڌ?'k�G�i)Y(�`� 2���o�|j֟.�W�X�vp����N:�e��]���_�&>�B���K�~u��+�$XZ����ܠ|��㗛��6�m�X߿{��ӺX%B��B�����Ӌl�4ӄ�e��Y���Of�uz�m&��UV-9��L<��9_׳�%;��������� �0�|:뫬���ZW�_躀ʸ�!8�=F�]���Z|^�������RLe�&�(R�,�Hte�g�WC�/vT��Ax�ԨΦY�dI*"�E!��K�>U�fM+���pߩ��j�r�1b ��񶫹Y� �G;�r��+] =PÙ(B���9��_L�$���tQ�yֻ���d\�����m��J�ӊ`�x@#E�v�fAv��v�#m]��2������\��'nX�)��x�z�� K����y�6g=�"�It�.�ܢ*�𔷎@�9���ao�h�j��'��4L�
��nAɥ��SQ�<Q������̛�f�f����	Q��+$���j�\2��=�����mU{ho\�ܪ���i��i��PbyJ{������aG��.&���nS��J+�B�ED;8#�Pv��DH��l7)�\��m��f8�%�
(h�2r�����K:�F���_F���b��46�W��R&.=�1cb1�W}.����8����4�ӍV&�0��\����;jJ�6�66V�8G�_\�^���)q�xh9��[� ���1���W�4��Z�QU�oy��8��A`�����H-�����Q������%�F)zE.�6{�����3SZ>�Ҫ���`
�:O�d@�|����-yVI�KN
I�r)��	�sR^S߭��t�2&j� _h89\��~�%�!ԗɌ��(V1�,=`�&�mپ�[���\J�6�:y�Ze��[�����ڛRn�,v�oʎ�\]e�-�	1�4��/������=z��E��0\��"y^��$�
��v��b3����X�m	���]�� �"cN7y�����qJ��ذ����ъ$T#��"^�۫�V~���5����U�,����?�a>4���z��#�I���U� )�+48�E=1Bp�Ӫv��"kIIv�Sn��s�O1�:��@��i�Ok�̛�~*��G�u�W���9g=���������ζ=� i.[g��N����d��h��'����cm��8��X�϶͢+��)xɳ�œ���]����l�%�mκ�h�^�|�ULTDgNk��/��D��q��	�孤K��|�}ԁ`>6�J��9�5�-T3���P�ؤ&Dc������7hβ
~ߙ��O^w�Bw��ۅ�F�L$���G"@��������וT�Iu�籷�1�V,�8�-��`�^G����WL}^~6��X,�Ӟ�0��av�䈔dyL��[	�����r�]���kE�7�d$dPN,��F�;0�΄�)�}\�q��Ky-b3�L� iA \b�Mjo<2�����0�mS�b4�>!=ݓ%����7^�-J�lrс4=n���L�"�<����W��hʉoL�Z�k�d#���_��A�=��y���52:�)JAs�E��z�<ܒ���ڌ�$\e��(�7�̷L>l0�7k�!"�7�F{M�dsmt
}��(�z͘���2��P`;�adn����}>�f�⚲g��$���Gz����r��b�҇&��"�N��f�ٸ?��x6��آ�:Fo����\�X���rx��,�k��2���2knh���g��K��y���u�{��7̵٨�y���N�_A�Gc���{�o�7�Њ�)T+,���G�4���(��j �w��+�y;A_.^�W�(P�t"� '�T�.��wT]ƪ �4.�f!�G��M����Z�m�_��'�}<;�ǂ�Ժy�g;)�\��zt�uYA'��΃��k�D�'7��'���FU/eGE��$p�H秥��ѠM�n\�_Bb 7}g��f��\it?G�<�?-��c��/U�>U Ӂ����D���8��EUS{;������M^�X�v{�J�`� ��&���>�"���S;OX5�e�x�u��d����V\h����5�=`V���r�i�G��~-�U��%����1�eņٿ�Z�_%&���7+Z?��uWm��,V�}�F��NR:
lZ���P�5��R^�c-u/w03�N��in��y;JJ��)do>q%_��e�м\��z/Tg���xa�|x~��;$�"K��%��B�n.��DRPXcl�69vY�j+&����ru��v.n�&���QD���Ye�11ü=~��;���N[�W���h<�x�� �w^ �@�έl$��}�iT���)��-V�Q�{Ь'�*���Zk\�^��ִ,v�W��{���åb�r���sU��aq���J��y7ҢLX�K����f�ZWʗs�ck+��Λ�4��':���x�2�.�:k�f�ͷ��c�*�T��D�<״z�m����$�*��Ơ�X��Sӓ�˗ E�(����`"������8�F����/�W��O�T(r�������(�x|h~�Ry��CZ;��-�~�hP���$�h���U�U��<���s�c[�.1�W��8O#���L��W���eM��<K���6v�,���k��|⁺S�0�E��Ŀ�s��-�
��sx�,i�H���J���N��	�#�8
�-���:Q�-;b@5fA����3�����P��縲}���-#p)�@�[VQ��g3����_���}�2�
�z�y�,�UY`c�h�hŉ���Xј��_��������%<K��C��`�S�h	�-w�q�s^�:�YZ�&�3Q��+F_�?8�l���!��ѫלڹ��>_x�v*�9��G�g7��K�p������h��YS����pq�{�JE���Zl���ꃪ,"�Җl�w�rݼ�?fIF7lUn�a��5�ȕ��K��^B.�)e=��7#�H�J��-�
뭢I�����5(g&�r�w�O�,5z>�~q)Ƽk3�#X���y�~MY����v�~�P�E��Os˓˲��gm�y~�?��&��%8�M-�+�?>XF7<v��1_fqS�Iz O��gw�e�Ie�^j��o|�Nt�ξ�oB
)�5u��7S� Bdd����#�W#���T�q�e��HX��þ3�Z��>bb3M���l��$�bQ����n!V )��z1�D"!��/+)"�mG�
,�g6=&����n������Q���]sU���tZ�K/._�%�(���� �@��|�:�	'Au�g%��.���F%�f���W�?����r��˛��0���J���m���oP�E&�Mo;6XX��@��,��*��[�y*���L�,r�n$�EO�:DOzf��B^yPG��zkB��[��/��}TI�y��N�?��0E � *�#��c+���G^��$�{jZ$��d!h��%�۾e���M�5��J��gxdo��g�����e�{ҽ)�̊*���a��\���j�
5��\� ���P�ל1=�R<) �3�륗�=E4�5��7�!m#��V��H3\�L���Ԏ�:��_<���JjbQ<��>��Kp[���_+嚳eQL��o�AO�,_\�+��hh�_PJλX�)=~�=;�R3���`���s)�薇�!g��^6_��ꪚ y�?hK�Г�؞U��YW����:C`7zr,/�r�s�������Vf��$���_����q�p�I�r-A	��ƙJ���R%c�c�yV�eg�5H�j<��kK*����Z��1�i������^�R�{��dJ&�,O��B�c��Ǉr�+�e�e[/��_�	M2�n����~����T����w����%o�s%Kʼ~�T@N��No�φ��v��z@~�we���9���}�4��{�kl�_�]�+�e�����ͿIM������0V�&��������𵟌�A�~��S�D㬍��^�7��2%?6�a�uu�}��wnvZ��?g�@*��ƃc>r��=6q��p�.�a�y�3$�j�+U���	@fb\K��d+�7S��S$&5\������y �u���� �<�M='Wծ>���ݦ��~߽��q���9������;����H��f]��M1���.CA�L/�m���>�����vc}�w#�hn�H���v$$�E�� ��Wg�n�k����=�O,���OH�Tz�W<��U�e��d��SRk��fL!s���Ob�&���Lk��K{|�K��{���`��%�$�C�������f��/�F����� j�nRw��t>�9^~�R[n�fFE���i<�77:KZퟎ�ݦ��b\�l�`t���pvL�K[#���e�������ˀf4�ŭRr�I{7p1��0xd�>��z��ۙmh��~��Th,:�V�7Fwf�m�$[�ΎT�p�A:�f���������������^��4r��v��~�q��_;��@��~��������Ӱ�+��u���{���!��!��T��<�|��<H��!I�1X��%|���F�C���6B7�C�rG 7G��ֶ��~����y�2��<8���Jn�V�y$V��<.� H�O:O��4��m��Y����(�q�|J�����z��^��c3uw膡.�H�F�e}�Z��׌�騧�����e��䊧�_�V�����Z��ɂBM3s�9�5��yv���f�I�,��mk���g��,=F��#�<5���3�V�䲮A!�t</*#|4!AG��Zz�S �{B��1���t�_�N�z�$��\�I��Έ��Hw8^�r�R�Fug�M�&tYn��<;ۊ,�>��z&kN��ZG�KܤW��3���t�3g��?�G�<*�'$��]���e��t!�z\vs����B��m�@����هټ$ݻ鐶���w{�*ݰ$�u{z�]�x5A�
	��ڜ`]�F��3���*��̟*ۗ�F�
 �'�Jo<��_;��Õݤ�k�K>������� ^C���H����?[��+�x��
��V���Ǿz��������u�p�佫����X��hC5K�/��Zf�`p�]�?SAҷ�H����R�[��"`��_�FՌ��ו����$A�����%���h	p�����%�6l?}���ο��\4a+�b�㰒Z�<<�'�	����O��z���K�1�a@�]y�ԅi�{ޝ��t�,63]s���rxJ�V�䴼*o2��Q���"��{�=�V�"-����V�e�3�{"1�ہ'F�Y2t}���s!g�Xm�*m�$�(��*�k���i��/;h��?�i�i�Q�U�5�o��O䬇&�.'y��I�6�y�ٸ��Ug�6nP}p�W{���-s�n�䔾-��Q ���=��$&>��#�k�����{���dݜ#�����/+|_l�ǷKR�MJX�Ahu���N�[?���!�_���b:W��Bw�5���o��(��}*���%^���V�j#�/�˿�Wq-_h�n�W[���"�n���q7��>qN�׉��P"^�DF����?DI�"�u���������R��	d���VF��>�I!f����������ÖCR[�+2æs֊�d����Kp�c;�td������QJj��r/��;�ȓ 7&rN�?��~X5'mBF�s��e�=��͜����{������iH���q��װ�D�RW�~^����� PK   J�X��t��"  �"  /   images/b09c32a2-0684-44ec-93cb-6718b830271d.png�"5݉PNG

   IHDR   d   o   %e�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  "WIDATx��}	t\ՙ����K*��mɖm��{��0mlІ@H����s脓�twfNc2��Y�I2K��m���p�N��t	��!$8L��`#۲�lY�b�R�o���ｪW������s]��=�z��_��Uq���G���^)�O�4c��(عs'.'9�v���'�������. �4� ��������<Xt y>��q�z/��~`a���b!ӂD&�	��Ӗ��2��`0�`U�'�"ԂR�w��R��Ԧ%I�N�RI���폞�~�(�`]�� ٥�Il#HL���M�\&YR'��:�u~���>k�Kk���1�����2���1Dǽ��t��t|�f������iig�E������$ 0�1RR� �oC�>B.����r:��,W1�߯��h��u%��<�S�|'�c��\�,�!w��}���~l۶� �QtβH���8���B�c��#t�Z0?���PI�P)w���>�X3�j�6��dH�&Ќz�!z���$��B�d�O%�z���q��a\n*��6�:��3Ϥ�>+W���z5�4�`zM���h@�
�P�!�!��IB�TXe����"�_m1cs����12�B04PkD@J��z��P�NAO�@��izh����P��Q�$�*6K� i���Z]��KJ�0��p���B����_�#[��~B˚�rͰd��dd?+:��)��;Ρ��3����S~��H%f>LW���1_F�m�6�=Q
~L�^�'�,Y���V����f�%я\��������a��gH��V�g�(+���x^��H\���,�d��%Cfl$Hy� �L�PA��:����D��0�ֳ�b�/��dg,y�~��ǿq||���d�&K]A	�|6bz߬Z�
��{/:::����~�y���ˡ�1�#�*�@2\曦�Bȅ�
�B*j�*�CtT���2GzjM7��LL�L%L$t�̘�M2��Qd�4(q�a�[;Q��54)�X8���(=1��ϠLMMa�޽x����g�K���[��ӟ�4ؗ׉��L��W7�UI?O�!���L�&�V"����`��TbVmDE� ���R�Ǣ�O �S$��y���gN*���~Ɍ���'2轐�ٱ�x��/8���n�2	S��'�П$��b]�]D�$tk~��Fq�]w����=�����~N@֬Y�x@0@Ӵ�s�,CUU��s|*��՚q(Ձ)#����yT� ��\7L�Ħ�׶���9L�~|d��y]3�2=j� B�l;�B��^U��L���>����F�$h���:�ı�	бA��G�Ʌ��%С{�KNfZ0��bc���CP|
I�?b~p���gOs�ҥ����o~�H$����'>�	p:��L,-###µ�������]K�W��c_�9���ZS��c����X1�#k[�X��
KH"��i�B�T��[j���
s�pm�����Ͻ�}e������ ����kjpv$��������Pu�R�Ǥ�U�����0䫅��w��.Ŝ����B�/[�LtX/�X�,_�;v��s�=w�^�mmmy7eIa�v��%n�Չ�EK�h�ᬼ�<J�vq�q�����3��|�l���*�o��:�C�>�$fdt���.�F)�p��!�Qr�� ��ϯJ����t4�H�i��3�_Q��%F|�)�?�/�D�V�C��>q.ˣ믿^t����<��[�l��~�3���\ �t�t�{��@�b1�w�}hok��GGQ���#T�#�̪"�76�����V�`ӊj��8�&�1�	@�`h0r��õ9�aK��,��@���8��,��>��n��^?9ImJH��o������A02�_�al��g�ο|c�_����o�ԩSx衇�q��,(��jjj��z������:�VS{��`�H~�S�Bmu�$b9���H�Y��`�V��2�[�]ſZ]#$b&m���H=���-�CH	a�f����#k;<*Ku��9@��"I��map��<�E�|hE~ztN� T�s�>{��h=����8�����g�y�O<�y���܎ͪ�;�l4+ �GV��ݷ����k����$b�0��
��rEW΁���*F��W�p����)�I��dF��)"�HF:+�m���pU��$�����J*Cu�( $� �N���,#T��M�ذ,�%I���R�����?�?���ѷ����t��c1�+��y�l��b �J{SG����֒�	У\�n�z�Uq6-3'�m��sa����E��dMi��f����J�Aɸ�a8.p	5�$%g� �A�����@H���g��>s%5�p��0��x��(��̐�b�F<*�0�7`�}&�9������n�8q7�pC��zQ�{SLG���m��t#��r�6�cܶ��/������SxO,I���Õ�K�,h�"酙��J�+%�<U�SW�2���n�f9O�F��I�� �'ia���b�6���GX���O�c��B�Ceb��������Cl�Cн`F�;F���lh@SM@H�4�q����th�5o�/$T�#uiݖ/(��,:�W:4V����M��E�����%O�%���߬-���$EKLb���8���a9T �CJ�QE�����.Ԃa�jʩ*����;66"�W�ў& f� l����^n�� ���ڀnd�(�ێɎ������M�����_¹�L(�p�x�'����9$g�L�\T <x�ֹ��I����`p��,�`k��1�4@�,�WBX*�Nz?��l��$���A�}9��	��g7�q.t�DT���Z���3�A(�ae_��/����"�/'�5/ l�2����v���a�NL�o���T���Q
�&�vro��K���1�َi��8�jʕ��F��]C���m�xb� NS�_()�յ��ί_ކR�hƼ��WL/ǠQ�"�"0�Ց[��u !�ȴ&R. �c�vaK@"���GM���VΝwS75a������O8n1rc8����Vzn���s���J�B25����Dݶ�^�y��HO�BM�zZ�`xIޞ�QU�'r��?�WK�<��	������}�C��L*�x���8V�&����C�B�V S+ŃI{!���!}�o__YUD�c���q��a]Y@x��Ξ`�`���5��� ���rPH�쌱H�`ۏ��,�\C\�Bt4ݎ1=YH�����%��|m-j������^��,��̩��,s~�Y�5-!ܳ~�;0����c4aDO�KdH�F*�B`{T��rdyKTH���q�^|Ј��6�shR.3�f�URW[W�p�B
{�"�g�lQ&�[[��&w�wxV@�E6��\B��n����V�`�@�@��A�%�+��v���дS5vZ����;�"{b���\��8��p?��K%�A%iXs;�+�d]\�Y�� YK�J�����I]�*j>b#ρ�k3lu���������J����3\4�®p}�6��G_.��, \�z��@�d.��O���^ϊ�ƒ� jC���v�j �%��(�Ĺ�0;�ɞ���(�������T�p�~�0��/̆�w��?��lx�s���o��6�!�54-;��J�5m12��9~5�/���IoV��䂌��֢{0)�r\�����іkk�=z|}�c�� ���3��)�Ѓ�*_2��&Y:V�D��T�EJ�j%.�3fVU�ΰ����ː�j���Q�vr��S��O�|��%�2��Mw��^���v-��|�F�vo�!^�֦��8�3-\5��q�:�����;�z�u58t&.�5��8q���F�쐦�����t2�W|�@�KE�˚"�d��FZ�̯f0�D��j����AI��`Ϭ�ڇ�K#��] %�p��R�?��9,���<�L:��1b�n|ܕ���h6ՅI:l�q���y�`�<U,�����~���c(�O��)��c��,�g#�Mm��P�Q6Q����-���+u��������0:��aJˁ J�4[B�ְW��֏�� �$)�/��l#�������A'�$Y��¡X������+`�H�(~ͩ��iv
7�q^o���	��؅��KG/0*���_�24c[�g������)"�z����]ᔣ�l��5�d5MsHΐ]�ܒ`���vY���iU�+�����+n���*���C>;��O{$"S�,��Ym$��Dqw����_U��"H[��<��\8���T�4qj��)m���?.':�;cO&�
@��篪:�>�&VS^�0�R}���Q��#���VS�P�
K	W�sU$'8���C��@�5zF��U��G0��������!�%n}� ���s +h����XF��
&
u*�R��W�[
UK�IX�*`�G�qeՔ�h\w�9���ޑ�=�0�Vq~�Nj����I�(ȥV^��96#WN�����S7��Rsġz'����z\���!b����+p�����9@��Re{�ʵ#������,!��U�A�<</�37�B9���s���B�(�cO,�dYn��*��������,���œ�
o	*���$�i%ɻ���aw�l���4�4褮�R�*4/yґ�Z� �	ဌ��3��X)	���+tQdZ9�y2pʉ���s?�)���
{qDQYᝐR����Ĝ�r r��DyPn������o��6�ХsOL�v�p�ݚ`;�G=�\_�,�p�f��ʺd�az�Gr�g�c��������:j�B�N^ɰ<`��f�3�!�[��$�x�"�N�Gg@6��e�ó���̦N��]�H�{�,���Aa%�ij1�j7��r��U�<��9�bu�"3b���1�z�Z�@���x�B���0�\}������y?�\���� @XJ|��")�H�,n�<��@Oh��C�±�s��z�]O�"M��}���Sn�Bnb��ΤtJ������t��{2��OuNe��*��%�;]A�"�MU��iMd}��'�b�"u�d#� ��,R�J�5�HW�'�H�Dɞ��4�H���(ًpIxGUT��@!@�Y7Hg}�H� �BOb�HAc���gr���q�֭��䋃7���J���b�dzƶ#�~q�86�m<=A�|h2#�֙�F�~{2�H�[��m�ھ)+��y��]4]R��*v�"�����B�U����d���
u�/
�U�����0�`��O�QU[�
�O��Y�ѳFש�ryۜt��nQ�� �>u��(�,�z����	�TF�#�;y�8�;���;����qj���QeF�����+��B@��M�$��V�I� �X��Pq���1�~RW�L޺�9`���9(�Bf�D`���? I�Q�*!�F� ����~��u��ho����*��@ΰӿ���k���	2E���_ !>��S�*�����XL�g��U&SI]��U=ˤ392E�'���H����p�7�0�?��������DnM�mi����%@�!���j/���W��Ł�I�]��9�u���>VW<W]�&�`T�&���E�r?�-�3��<92���Q�[�41��I�p��f��!�59�oy]`���~������~����TY��P��W )A�����VSܪB
�N�U�8wU �p�e�p� ��֖�Ʊ_���������k)^;_ߍ���s*䳫��ZE�*�1p�ݩ����%j���殝Kk�*9�#X����;�eU�2=K��-+2��д���{ȕ�׶�X:�8>.�=q�#9QZ|l���o�j\��M�f�䵯\��[&��������
X�M�L�jQ�U�J\�+��2�^���dZ��W:���~���]O���/�d�Ur��C�"��VB��WJ�;���B��]�V)�FN:�Aۣ����O��E<or�Y�c��1��y���(�U�� �V�0�#� E)/�H $fEck�U��g��}�d� �OO��h�T�R$�;���LR,ӄ�� ����TO"֬a�)	>)_Xu�-��Ī�������ª*F`TS���08�����lF7;�Nٔ����gz�#nP̷Y�HIt���1�!NAMQF����3C��Wmϩ�j�
^�.����]�FE����
x���e�=85G%Ϭ���jM�ni��bW� �GSx]i�к�U�_�6P؈׆U,"08����QL&�\���L(X8�:eZ�v6�s�fJ�P�$N���5�O�g��'�	�b��WMq6�D�����*��7����He��F4.��T��Fq����gV�$v�{�8.ě0�����^��M		���i�4d0x��E�'pr ��<���c>
�k![sHӼ�lY�":�'_�l%{,2F">�0!�hZڔ���������HM5T�t���;��YD߮dp�A`&��wP�y��8�<���],�o��x�[�X�YX(��Z�`�%���=�;�*h���NM�{��P� HN���{!�8������Wan�3̲�j����QJu�_��,A�����}��H��#Z�[x٧D4Ͽ���c,��* �M�}d3��p�����0E�Ob`Ϸ]�Q�.Be��!��Ǟ��8�@�+��������p�r%�)�d�D���Ŧ{���O
5e��+�9F0��9t?�uq��>����8p@��H$��o�^T�Aihm�(��]a*��sQ��*ZHM�O�p�̔X�D�،B0��"�����}�wsm���C�8�Y�~=^x��a"o6�ڟ�����$(�>U�
ט�� �J���4�^P �g&�?�L��,`z]��0�Y;�۝3���`^��͚��q�m��G?�����������H r��� ����]P'G'(<�����Pm�;K���j 5O�q�����Z�Ie� u��C8���8��d/���y��w.M1+ ��WJxSĻ�gΜ{��w61�����C՚O�E�VqO;'k� ���:DcQ��0v�a'e�p��NabF#�s��$偢�>���O�����ݏ7�d�y7�t7���f��ɓy3�����<���ػwo���[OA�>�؍��q��'7��5^�����XԸ���A"k�>b��"<��C�3��ΈAr���ǜ�%0��z������o�����g>#x�+w����Y�cV@x7㞞�k��0ߘu��?�y�x�ؽ{7z{{ņ�_PDG�֝�GľK��+u�(Se/����XD��L�M��&���;s�N��Hj"�(@H�j�"�&���{_��#����#hoo�֭[��p�j��{�<x��$�E���.~��<�]۲a��[�Nܜ�����������7�B� h"�R��p�Xb��IQ��� ZE(��J�禈�~3 y�C���Ѡ�3H�5��:j���F�(KR����߇�����{0��C<'o�̻l�����2���b��hN��%��'�ă>(����5H�VUU��`�{��;Z�Qîs�8;j�$����R"�2����\D���-H �w&{F�. wkbz�A6�tV�[Op�y���HO�`0�ql��M3l�յ��I����
�CCCx���199y�0:t������>���N�B�y|j���kh�⭉F��'u�A&���%��[���F5� wҧ
	b`��c	�`ˍ���w�;�&&�R��<]&g�~���!� ��Gg�,j�`n�ga���o���w۞��
ϝ;��{L�oK�.�Rq_Vxx����ͨYy+tCE:1C=U��2]���Jf`WNrc�V�4/���ܼ��:�%��I{��v]Y���1��{�����������bO���r�p�d��P��Yr�4�	�FӇ@u�-0I��4S��5��9����8�㽀� ��<��缠\�@��$<��W����)\
��"�S�,5^>�R���uk׮�jvf����(y`zÇћi�D�l�L�,+5%��<p�
@9���z=���Q9�%�iH�´�~kyKҦ�+���.�濉�2��2^x� ���w��7n۶�����H\�Zx��|���j�i��ѧ7aH�!�˶�/�x�j18%��\�H����!)�:i��8�F\��������[쯓��7�����{ǻ��p9鲭�я~�=���W(�!���9���G��L���Y���2͛	�������3q\�"pr��d�[,�_�$��0�0��"�U�E����DF9Dl|�Ν����.���Q�x��$⊙~F����B�xj����D��f�6ПE�a�ژ	��&y�w/�?F��H�}[���M� ���L--�){f�d�Q~��?���lO�@!�8B����4�5F�Ӫ��	�F£�*Fa [9���$a1J��İ��#��x��Aa�V��X}ir`��h� ���"��˝�����r�IEMc����%q��|����p�-xe#
V9�t0��0Y����ZP�xi�#�˺�ge����xj�|��G�B�H�T W]�|Ш����hJv�)�    IEND�B`�PK   J�Xr�>�� � /   images/b24f041f-17b3-48b1-9f28-cb1f31b050cc.png�gTSk������H�o)қ�4K�
* UB0��A�J(�E�RUB'�P�I�ރ&�jh!��Z�����1��{~|�Xo����|IB訝?�v�����}�m%g̟��'�_~���p����O����s������\�����Mv�􁇬n����m���\���p������ճ��b�.��k�lTTQ�Cn?�LY�rp���M֝�VOY��u���h�~f�����y��$+e�%+��2I)��ywK�*����ƋAg�?��+t^.7�.p&��NG��wg���~I$�_��i�"�pw�e��͈�t���47w��x�[��� K��ӓ6������Pu��ʏ�/���Aa訨,��x��
3�Q�A�4�ɉ�U�5F�0`}��{:p��$�]��I�ץ"��' 5�x�!�A=���=����_�L�M�Jj��*&)�~4�Y{�o������ }@b��D���!��/�+�M��u�5!�;,Fə�@7��jv.���ɛ�++=w�-Gx6�Ǎ�'���HQNS��:����>�gE�3���Q�Dha���^�-0�[��U�����/�a7�Z�|��d佉	��޷AL ������&�`HU�9���?n�}��!_d�Y�9Ҭ�	s
<�w�Ԕt�h���Ip?���T��.���ͽ�W�:h��Ճ�P��X��o�N�^��n-Nդ{�b�/4�՟��σ���zG��`�����%�&���oX%Y�*�!)��#��J&������s¢zG4���%��(}�����GY"�G2Uץ<
Y�H�Gh4��'j��J����6�7]��	�&�!ٱ���u�����Fc�4i��4=�1Z=�0�޸�/�X�X� @�F�����Z�W�q�8��ya>pO�7R+�Щ`cc�ű��8ȹ!7�ly�<)'iQid�LRc���NaUa�7�Lړ�����#N�U/dX5M� ��5poO,��w����5o=3�奚��mm�U}4),��Y_���ܳ�ߢ�"dе�F:���㴊�z�F��U�E�0t{&����D4���M ����J�;���x�ϑ���]5SJ�7���a0�Jvc15=�or�}ʅ�Zٻ,�*���}:�Ѐk�^��~:U!�1���W�Y��cuV�`�J8^�m9���@����tЛ���8q�v��7+��8�����)2UH��P��@vE�v�Л��{��}	�%0f�H�"�9? �L����{6����n�?g�\�:�1�#�{Dt�f����g�����pI�t"��۽���d�9��H1��`F�ܪ�迫���>�E_�y�5���tz^����s>5�5�q�^�0߬n�u��k}q�*��[��к���,(�7�JɌ�V^x��a��^��MW�Pt��R��l���Z��,���e�-�I��M0�.�����۫,�c&��*�C�9G�M�;��v@(g�rw�5^9���7�҉��H$RRq:�MHF��c�?���Hy�f�X{�<�!�;��g����\z�nvj�s�ժ��*%��0��+��I�������z=F#33�����Z:�#��*�x
>]�0�������C���<g��6D�1G��f]�$��>�����K}�|��v%��O��:��L�|��r
DĤnԎ��ld�Y��맑{�����ޔ�T���Z�v��
�����2�̶�ݨqFάP�ԧY�=�܄<�|')1T�!R>���{�����0�;����K�V�����<����	rq_=]�*����n���*'=�Pg ���g�~v!�y2b=퀕.?v�ui"@P4h�z�|�j�Y�u`�xvx����<��e��GLpo��n����5���V�ꢃ:�5�U�H����O�UN:�O�_���~�)&��Cؗ��&N��.��RsQ �oe�^����h'5}�k���?AC�!���a���'n��i(D��*���H��Q^^���x��qu}w�����O[�Fsz��ir��&�/%����x-q�.��D��!�,���@���= ��|ډ�f�I�׬h�)ĂUI�\K`%�*�1?=�UL}���4\ͅ �~��N�����x@ !��)���}N��z>�e7��>D��19H��md�+����8�ſ`�A�#��#��{�CY��/���!b����[wÂ{
�,�"���د˛�dQ��x�����0�*�t挃t隒o.R ��"�WQ^�6��6���u~L��4���:V�B|KP�����55�7�#�aQ�}]ԇ#�kY=��q�R�����Fh��❷j#C7kF�, U��$�_4S�������wF����ۋ���4�G�iq�:󪲊ѽ>6h{�eF��V�XA?�^�c���^��Cʁ�F�.x� ?Yc5��2�V��C_����7�`�RX���(���Qz�����d�7�)q��S�4���GARzz:��+�����#�j���몚�%Y����a�I��*�`��1\�Y�>�Q�IM�:�U"��Bkٱ���.X��bow� �������������� 2�|��=�B�ƹ��wU�k�~�����x�������_��B��H�A�r��¹��P�%
�a�S���NN���`e
�4b���AJ����eI#,�q�;��������<�(��b#�[g��v&n���j*S��	���
;��V�ubM���w��Mi�l�2YW�:�Sc	�����~�i�}�����xN��U��ѺQ�c�mV�%�4���ƪ~=���@"�I�/Q}����
M���x�2ɡp9)
��9����TĻ�:)��(�$�W��Daa��+�M�A�	ѳ �~���ď�
�"WC�3�z��G���{��@T̷�~���}��6����JPu�C�Nܛ w0�76�:�`?�Z��x;�Ta�W���"8�#��ȉ�)D�<��uO�u���c�B�u��%���XOJʖF�g,�������*%b��>��N/��������N��HM�WA�4��M�n�H�˫��U��#%��=(>��`j�S�Dd�]4\�K;����U4J/� �6�# ��x�{ͧ�ۋ�<v�����n����vuu�ۭ^�w��v�ᴗgu#t��l؛���fұ��$~�1�ytMC��p��M�ܴտAx-��{�i��8ֵ���������B䳣G����߳�(�; �!Fft� .?��Λ5Ҕx<�y;k|s���&^R$IQ���"�������zz��"h,sn.�C)�d�����H��O��X�0 N	)=�%��d�B5?w�Y6+�N�3��I��2c�q�05Ymԭ�F�!lOR������W@�X�t�Ͷ���ۥ�U�R�X�-���B�OVL���6��ᨆ�
le<K��ӳ\�����_ZZ�RϢ�F��ue���B�<��Y���'��{QB�\��&}�Z�oա�Ǽ`�Xz���P�KZ��@�/�4S�����3azn��sd��MFg*aYD�pZ�eP���}��97��t���y5J.3߬J�P1*�k����t�0�Fadg�k�z՚}1�=tӽ�5�v��<���/�0�DH\h���ù+����*u��u� �v�	��X(=�G=�x�<�U�F�2Hu�l�L�O�{A^��@�'�i;��^���9���t�&=�cK��� W����N{���,�~���J�G��!�C���E��׵Y Vw����z������ĎVY�79�'����k6�_7,f�M�"���u�<oM����$�<�.2��Ë�l�(��J�̯��@j@5�H�DO��[���sp������_ �(z�� �?����]�=;�p��un)a:ƭj��d晴��W��̃�����R�r{�\=$qa�ȿ/�~d9�%i���6����ON�",-�<�&��ڬr�mU�7Ψ9Ց��׏�I��X���ǻ�޹�KJ�K�X�5��2 d�J��!�
F��a�moDs�*Eێz�~mL�/��w׌?����ܱ��t��1����!%�As�����5l�j��f��ڬ��>��ƌN�Ƌ�n�&bJ����W�3��[7��Q��:J��\o�-�����,5ܿ�D�m�G�Hሂ�&����I��G����(��X]�C�Y��FM��ВIzzc{�j#?	�ze�u|�{���2n5�CaZ	�*���uϞ��m;u��Vf���[!j6g\ax��1f���J bwR��iF�&��f�pd	(���a���?�.��_�Ά����{f`v�Q�3��Ī?���>Y�"�;�h!����4�}/9L(�-WHs�O�b�8���]� ��u0n�-o����g��oZ�J��x[@�i�ajJZEO��0�:�b#�����dL��Uި��"m�?#�<W��`Y�����՝��}�0x*/�ͻ�2]d�Z[C�c�/�Q#����W86�]��:�N��L۸�w^����f �7iʃ5 �.���쳳>�L&�E)���O�x��̥%R��c�N)��!d�kۛ��P�?�pt ��+G���L!��c?�U�M)Z�>�K"��@[^g#���X�iM]*k]��DD�,�ظ��!��WVt\>�I#���[�2�?+���u
}
o8<�[��S��>����m'"@�g�K.�1����B����I$���RY�|�f\᭸X7�:��WFa��(���]:�� j?���~�����G��e��^"Ϥ��? ������y2z����M�ˢ�+j��Q$ٓ�ha��b(1M��Q]�I�t;$$=�NQ�~�Z�FW��� "��QS���N�Jð�l�%�*�X)~�*�q�W����ܙ�O�q�D�$-��N�5q��dk��oV�������Y� ��|���
��G��6�!im�+;;�t���*F�="$����"��̠��6����ƶ��ĥ�ɧ�t�n� ���VR|����������J�Ϲf]�X����G���C;�G%����?�;K��O?��6|dy4���r3g�;>��f�2����$J�zՒ�M�d�-d�q��.�����!�lYi��=}��{`��v��v��(�����H;J���'<556W5����{si��駕Fn���&��/'��u��5	-�F·������?�g��`�_�g-�;�	��H��U���Q ��^5ЩE�
��/.�o����'9����>d�א�vr*�}%l���I��@�zP�rD~J37��):a����@fr��e����������w������?䖿�� ����m0��J�a4L<y�)M��qc���_'2��[�5������>	�]��j�޹P�쨙�s!�_�F�W�s.�|�����?�]v�{D�x!�N��H�)�DKK{�^�&n*N���h�=���$�g�|��ύ)7�.�������{��yQ�nY�eJ�P�TP��.U�U�g�W@K�z��z_����w܋�͛?͛��̤�[��3hzr��U�L2z9�[�Ϗ���as���Aq"�`�q��>6u>u��#5�
�2X�O��>����h�*�*�W��߻�P贆݋I�C?z�fL��X�sC}Sna��to8�8+Xɽ�A��\En�ʄ0f�gG�B���U_z<aȠ��cPs3DƮ�5�h�r�}E�{�	�ꎿޓ4�U��j���=�������?rZ�a���ѭs���iV�W�����lFDN��W
H}>��\a���`��=�I	7�x`w��_��U������뵳2L������'�+�w\�٪T�e����[����W�z��;��"�VE4%FDb��?iѮ��xC*��g��z�h�]�pn0��=o���i�{��U7�TQqq|�LJ��۽�K-ǮV���ry���o��+�u��h�D{���?���7�zo�h�j��x_�_�ϵt����~Th��Z�����ͣj��="v�H��Tq��z��k漪�<�����b4��
�w����f>h��֫~5Ȍ��g[lg�0���WOnn�>u�̵�h?x��j�o��*�C7u�f�T4xc'��/5SvcĹ�Z_�%�L������A-����,_kn�_�e�O���L�^���"�{�S\bmv��h�1͹�� �~�v���3�i1�'���l��l~z����.�nM�u��J�G@��ݏMO|���H�f�+8|�^[���K,���ӡk���1���_ھ_�!`X�.�Fh6,�(dG�G"Hx�ұ�9����C���+;+��O�""L������"z`ߎ�E�`_U���^"������u̼�B�#���鿎m�u�.[�8q@}�:=���whb�N��V7?�ɣ��N?{p�������
��(t=a��m�3�/L��}��V��(�s��"}�^�ıe����՚�PU|�ޙ��1��t���0����9��ζ����Tc=!�?Y7m�g�R�>>��fڨ���6e���r�8An3��N{�̝חr=�_yȽ�	��q��\�t���r��1+�8Ё��(��+������,a�{�X���\զ��ߎ5�8>�R�c��1���N�I��N�Ѫ<MN���D���8��.�����Шf��ǥęF�G/�!�<�̹�ǬK�6����y�
�Dպ�r�:ҍثs�֨|:��ZT�}2��-�B_ZF������Y��6!�ֹf��|g{m{fǼ����kRaN�"�n�T���f}��KZF��ֺ�����dW�����+M�)�{cm�T�7�wj�E��a?pVb߸K6
�%���u�;�u�~�Z�����-$ۉL�
7;��������u�#�g�Z9VLnt�a��+֣�T�G�s�b��c��hר��ԚZ�h�g�yç�}OU8�W�[8ȁݮZyY�e}������ރ5�V��j������U�q
�'$k�{|��N8���� N�d�����{N���z���V*�3&��j���h"QypȀ�)�]���1�l��?��{��ɤ�W�*�\U1������H�}^��XO�b�A;*��vY�V�?Z˭�fԤ���;����:I���Ѧ���V���CޫIF�ǙO�Lt]��\�
�_���a��5��Eu>��k�
ǚ��3Bj�>θ���>���J�~ϩ����k
��=L�șઝo�ǔ��|��򆖧*T|�K�Z���E}t�q�t[֮pZ_^4��'q���0��Y����G	)�
i��f��}��}��{�#��F��xb���1J�t�S+�� �{��'�h�]���������+B�t���H��`T�0����b3t\8��O����K҄�4���kw�zjD�qV�hlLsVk�Wt[~_1�B����'Zm�ȯ��;3M���y,u�yV_���8{�`���k1�Gg����ś�+�z9�ʍ�o�0�s6�N�7�ä%�z���5�BMw������r�Q��iP��\��S�q��2�� �C���Z���@��s5��aڡM����,���#�+�'�׊��:$',�?^�>ܪ���9w{���d��=���q�6����o���8�����i���U��{$�'���e��\/#{����1L��m��ð�q4S�~9ͩ[3�c092P!����ʵ7[xv-�y�Dc��k�Q�mV�3O�v��������-&��Yу ղK�����)��)��/?�z�*�щ	�_L���o������s�E\�I��ڒ8�r?�uB��XF�����J�Y�����6�te_�\�v�}5i�ت�3�YJs�p5��v51���Ho��=&	������N����,ګ�>��-v�w�T}�=)mڔ�>�$t@Ajw5-��y�|��HX�F�f����=��%n� ��z���4��[���s/-j���c�͌	��ֺm�M�F5�����g૓�/��w��n�E����WS���c����p\�S�ً�t<�/o:*��=&��v�>J���(}�b�pE���s��B�GH�Xo��l1�Kիxyy��n3�^��E�����c��_�s���N���ʹ_�.��W�Z����K�c�}]���\P�}/Z�k+�Ć
�_9�fvE]��wT�$�91ϰٍo��kj��s���<�vb��e*�&�=W�1ȟ���]-<�Ү͎�2 �Ē�5ym�Ѫo�1����_$]��c;#;?���c#6�rsp�k��i�4�-�ɵ�I��G�k�����1d�{V{5Y-k�
�`��<��)�mr�I�~Q�Be^�9�9:/�(> #*�p�p�<֋�\{eS���S�7lO'� z|�~����>3.�&"�q}6�x}���lpr��+�ڐ����Ne�U]:���gm����oNhVU�f���A���%��;>����䙵m���ck��]���S��?�Ty�漏ɷ���0��8@M�`�N��@ ��G�����{
H�9�h>KM6oV�賀����^c�����>�>a+�L|Bqр��$�������:�ɕ~uִ��9�Rآ����}�`��q���<��^K�ȴ�B��Tb7;�8�k�]'�%+��]��%�������wT�T\�'�e��L���E�J�4GD��phX����#�z �qn�{;�)qz�}�C
h=�Ɍm-)�v�Pr)��V�鑎Q���$��ȽRcG�x�枛��������k�4^�{�ve��|�_�'���"J���xj��F}^�CqV)}�M��rԛmL\ov�^�)N$���Vu����L��D��F��͜
�05]�r�����K(��|�υ���F��=�"�3��%��hi�8�ū��n���kKUp���P����ܣ�}G��.A���"�e�(,W�K� �����H�~�N�:�����S���Ee;��l��F�I�4�WO�y">��	��$| TF��yYe)�2�0т6$~3�]�I�յE��Z�o�~S��sũ��"���	���G�/W�p��}j�H��}m��~�Q�i�x/"��j�䨯e�Ϭ�.���)%F:����rk��֬�&��r���m�ĂP"h^�e�?�f}�|� L���M4Oymg
**�l�;�V�L����IeqZp�gX��%�l��)��47��}i�����4�,�S���>i�>m�>e��-���$���*D�hAk��g+��rh
�m��~d��M��rѕ�j�5�����L�55Uj�/n��P�%�\X׉�Ѳ6��'��/%NY�������E��=�~�`iڢww����L��W�|�B�j�_OR\1�P��G�����?�>�?����Q%3�S�2NB{���!��4q��Rо��[�3R:g�<�_�P%�~��������������b�~RK������A6��iD޺W�/�r�ѿ��%�F�W��3`��3�y�ݯՋ+1�
Sу�꓿n)��H��
չB����BS <��q�J������M����K��l4����I3h	��re״b�X�ۼ��ü�3�tU�ա=�,&/�з��.:��b���f���ѾA2aS)h�s ���C�J���Bű&��ا���"T�2A	
��i�-�4�-���zJ>_����m���9��'L���8��@�^��xk�i(% m���V�=b��jٲ�%�D-q��Ep���g������f5�Z��ĳL ^_�<|����,s.�R����Q�%;z����aht����ě�E[���5�K�K�W�s<���!r>�s���GV����o�]�v��fwC4{��\�w� cH��X ���Ĳ�Am8�{�<�(ThU���ڰ�����˭���7�;�r�x቎�%�Ez�����*vU���'Zv���aw�Gp���^ʆ�O��k����^�<��
T�D�_V�S�~}���{����)�j����K�:7M�1�5m �P�&��-�`�ok��rv~�"�!?��h�l�:���B8�­�/ʤҪ'��լ_�i	P��8���D�%Gb�L�&OZq-4?��3M��V��t�K����cW�E�
"ӗsiH޹ɶv�H�˱��c��^bɞ5iw$=o5R޼=��"{�bIa��*
�29���x#?2�(��;� "�t�M�nĈ(N����$������Uΰ���Qx� �f߿�oh7�V1ov����G�!��Ŗm)0�fS�E(�E�.Gp"�5��=;m4ڇ�c(Tq�s��t1�2���R������Ae|����ĭ�~��ms?p\���Ӱ�4V˛oq�r	����u�>Bˆ�~ey��k7}��7��0��@(��ߌLA�pf�?���2< o�P��gB��P�[�Io>������d��c0�̵�H{㸟��Q�W�n�_���e�n�5�5�9��Diw!��9R��SMM�ԣ��X>znfn���|�d�;Ϩt� �v3��n{ad�ɽ���.B���4�-,,�)}�}�V����R���G��&�Xz���-r}ru��"�2�����O�C*#�ڿ�S� � ����.�LS?�|�fzc��W��pe�]n��m�4OJ#��P&��ֺ��%?�����^����dKtNSIȂq��m4+#&oχu���C~��i�@��oF���|a�4���'ٷ�L��.�pf˘�mݯ��Y��u�7��b�s��.�'wYsp�(3&��)@1ނ���T2��P�C�̧�:˨����.ny?	������aϣ
c<��w��R�2����m��m��)O�����~X?G����]�#��+�|���%��������e�����}����o���[���ږ#X#tP��+ƫ�M�KmF]u�M������&z
8��&��6�]y黓�R{L��<.:�PM**]ˁP�ڽ؏�vC���r;�|C-�5o8�u��Z[|!��w��� ��ڧl�'�5���$�d��o�S�� 3ŝ�[��Ͳ�n�'�~Aj5NR�ʂ�x�<HA���W� ȧQ��]�w1^���IX�G�7��0Xզ��n��~󼖘:a_�
�Q�/W$���'�T�*�`T��x���u�g���͋p�:�߭.��Ŏj�����Sh��ҷ��e5�y�)��:�0n3)�O�
	_��J$�(�Z��_�����$LXd�$��5;�R0X c��m�&�23�7p�P� ʦ����e���"V���?��%�V б�L���5K��^�Z�ȕw���s�NRy�5A/�`�̭{�"fХ�H�v��ﯥ�J�j�9��r+9�7�ŒR~zN7=�C�,f 9򞻬%}��x+ܓ��D��65U���f�r���oxC�8�> �NE&�t�	#�<��|�g��X_/�ޣ5�M��	r�G�#vc.��ME�%ht��_�2-��N��|�Ԙ���\�,�:���Nl	-@�p�S��R��v	�
��� EF��� ���<�
����n�3E����WH��'ld���.#m���x�}�J<<��؂�O�/K�~jy����tP�_;0���L	���b@7����Ylӕ��<]���iSa�:V~���u��^�*��4א��B=�y�q���]9a@�F�в��{eܕ���%�7!2��J�:=�h�/_��D���u��x�h���G߈��Dו����N�Xo���(U�|f��VK &�7��%�IcN$͗K�p���x�"G�JO�v�s���Ş=K��Ƽ	\�sY�-���>����U\�;���,)JM�a��`��
xg����u�\~ $&��+.2��n�O4i��#4Ǭ!Y� |����7Z��d�3*6��!�o,�.���̕�� ����#Ϸ����̕bC����<0��6	��h�~�吻�/ۙ��I. �5��ȂzB�!�ky	��L���珺�@�V���I�#�B�3�_-����,>�?�������g6�zV�D��p��'�l�3hj��]k�T��i�W�4e�n�m~��|�Q��2���T�S�]~jX׫!T&���P��[�3��8]xk9'	�&(Z�m��0k�P�ԩ��o8��⫑��#��1�N��/�KT>��@7��#�)[)>�8#v�$�L���DPl�	�d?MEY����6�q���i|kԫJ�s	o��B��?'Fz�|u�x[[�Jh�9�
��oM���DT�� ��5��=��7���\��Xjm�.G���H�.�Z� ��#��)��	���z��1<N��hN���m*k��>yZ�P3:�wܦ�ޱ����͠º�}n��	]>pb%	�`�w��@ܝ��~��~�
֛Y�G���P���̳Q8�+��s�8�o�$v<=kW�9�Q~���b�n�x����Q^ z8Ʈ_/덈�.��u��N#�gxK����Ӌ��������ȷ�x� �d����ӿ�m��%�|��n'�qyK�h��A�n|Y?̜);��L�tX#��%8H)�W%L�fyS'P�s�odQ�|�eD+A*�ۀ=�[�������y��Z��}�������vD���� �� ���Xw�@Bޱ�p�����s�&'�._�B�&72LEZ�Vs���*�"�?B [ n�F��
4a �c��Л������?.��wj����Wc�;�Ŗ��r~\P̶�n~[>V���cR�I��R���� ;zPa����i,�.M�"���s��}4�x�)F��g��*Z�)u���);�E�r�kG�ͳ���Y&d���� �[(�������6�X@8M��ID��9'M"��+��G�s�H�9���s+��;눏o�[�� ���7G��*H��7l7d�S�y�����_�����*��vw;[=�(eNT����#y	+@����7O�� �� �����"T:�f`��Ҩ�2�ĨC*�N�0�/�kC��kna����D�Ȕ��d:",��z$6��'�t�q]�Kp�F:�j�(�:xd��v,tQ��f#�G�Z�k-$4��X�b���Z��daO����sT;FB	a1�^$ԣ'$����G�r�.b�v��mQe�ơ�e�<󏾻�S���Q��m�*/��J�4
�@%�3Y0|�O�T��5Tf�?�\�C����Z�"��ݩ�U�2;�	����s����ui�{:�Z���ɕ\��ʅ���u�-�
�����y�LMx+@�l8�=�E�Mx����Fj�j�����h����w����@��3���S�6T�@53���p��2�*y���K+�ۓ�*KH�$�@�0�)S�1����X��~*�	n�˪�{]��Q�9t.�g�V[�0��������j��۰7�O��\A�UPg�=_^�3��j�hDl$N��k���f��>�8
 Y�fZ���` `��I��t��0uўzr0i3�5��Y[*���>(�0�-���0�q"i��=|�Pц4#3��nW��c���gJ�L2;��\�I���P�>�y(Lƺ������V�qSۻ��0�a�`�r}�(#� Ʋs���g5p��k@l����g��X�n�"fٓ�'_���0���}M%�s[�y�����j��Թ���2R;�S4�{��HTlĨOΞx���Yx��6w�Z@t�Dv�aQT+)=���i֓�pC�%����8����D�����	b&\�=�l�U�ð@uܷ��uM@h�ܽ�Ǹ%M��g�����s^�@�mZ�_�yY.7�5lݼ�q����	��Y��M3;s�'�d�FN�/��s�ܢ7�T�A9O}�&
���\�@]�d7��bsR��w�9�C��&i�݇O��.4���VH��L2T�~ �fY��\�2���L�&�R=fL$��_��|��w�-�ԡ�(�������v��Q7��`�5́L3߅�@�f`�1&^�#S�x�w���a4��m�	�{�����<K��Xw��מsR%&��7�w%��u:�tXF?wn�Sҍ�J�aC70�A��͆f�hDE�<�����G���|�/~SI�E�l�U�K�u�*q��m�>*� ����CQbu��u�I3�C#�N`F��Љ����Dm�sм��( ����~ �o(����W*���\X�t2���4�tQ���kb��6gl�Z ������[h�*���_�H�Du�e�&�% 	�:��w���M��~��OԏtƔ˙���_��x���]� ��=�@̱�hȄP�t���5�I��{],@�����U�q�k�`k���G��Tx>u���R�+��R�.��l�����EB�?17j����om^kdRI�T�k0fQ0��5>���@yl��e�1�V���1")����v��K�h'���TW�|ŐG�w�XΩ�`ϑ�2�j�?�JMx5�
=Ӷvʭ\:�N:������g�|�7�H ޴n�u8�p���7x]� �^# �l`�^���;(���o��'�Or���%���pVj�-~�m�7h�{��M|�1|Rh�R[��`xi�L�Ӡ�4hC�=2�F������֐�֜�~avi�d`G� ��H!x�$g>���>�唋�
s�/���
��djMQMؓ���&��9�lfi	9�����DKrݜk��]ǥ*�0��ubhw�E	�i���*�p�&K`X�3PI,"=��?C��dŌˤnn�ܣ(t
n�� ���aKm5 4�q]jW��K�aM�|�1�7  ZPF ��|~��5g̻WB��P�����}�≘���O|F\_Z'�Y��:�(�a,"ah�5	;�������_��� C*ҭ�`#��$���?�c�[��R!~�hS>�=���M�f�����(�	[�z�/��dL:���� U�g�|e�`�ª��(W=�Ђ�r�둎4 �����/VuA���Z0��U��P��J��Ե�@P��砡>e��W�T���tZݫ����z��Q��I'�=�I.�ɋ�Ϝ�RNh�]��;�����P��g��l��������3��7¸M��l�#��eE��^H����!M���'s>��6,v��uߢDE����O a.
-��'sR�M�Ō�x�i[P��|�G�e�b�tC��4B�&~䪗r/�pR[�q���]�[?�bƕ<�$��+���5��:�Dy
��w-�֛K\t�������s��:�ˡ��w%j��?�!�s��G���ں/I�Z�`%��0�f5^L�LhG�f�f5�� �o�y����j�A��4h���x	Y� =F�2���q$��hK�>T;I (dsN�3C{M���%� $O7m�{��2������p�S�4C���J�	��Az�!�+��Ǯ>ZA��kBk�p`�@���La��T`�r�L�qC��@�rĔ=���QVd��׊����G+ �<Ǿ�۝��;������JLK�`X�j�= �h�(�d�{�@��s��#/O! 9ۡ����C�r�l�_<�����g�0z�&]�l�Ǆ� �%�7Y|+.�T!�TU����~����NL\6_<Zu|�R���r�r�_�퀷_֓�'�z�2׶�V�1��L�U.7\��������b[�tȅi����sL�;G�u,|ɢv�2{U�vOL�e�<���$_�}��U�%�C/@��� 5�2��ÇOⳅ�#b��^S%�
?L�o�h|��A�Y<4�,,XUU���m	���04�5��c�Ix��|�\׸*/Mw	�5ι~c�|o�� )��·��)F�&����o�+:fїO����w̢{$��ZR
B��[���+ܯ|�t��ظ�m⽃#��J�	�͒����و��j]b�	�"�5�N�G	nu�������v�<����D���]�����*6�]�70�|��W_a�w8_�����(���V]��ݩS����nvdI$�|���m/M�E�o��y���t���}����J��0��[6)�{`ĸ��0-��F7?>����c�ASQY����3z'�{�3V���#��^�8lk5�7gh���{AE�����V��8b�K'ݓ�����{]w����T>�#��L:�
¿�U����4gO�$V�8�\"dciJ#N華;��ӕ߹�T��;$�Tn�i��ԗ�l���9Κ�gۜ����|Y�1�C��h�^�S�4�dU�C����ۊ���%���m����@��7 ������X5�)^��#t�1�B{ř�D���g�V��3��l=Zc��'����ԕJm��N��m�U��u�=�tAo��g��_Eq�H�gX�����j��tu����8�ؓi�=2��%�;���t�z>e:5�n�L�Y����j��*�5�RL�3�ڟ����g���|={������%_�r��j�	�M�x&s��}pM�ʧ�֕Q�=��˳�\�x十͏�rW�',,����U
�̳AG�OU7ߟ�u�]��b��<2��E,��l'�lf���췌�n��F���ò�y%L�&�H�e�3�OT�i*)�������'�f��o�G��߅V��H	�O��t�sa�FfN�fZ6�ę���J�=G�q[ �s����)|)��]��K ��S�<�W�؝u@��N݅����m�%��ʱ�4c�^�[Zh[g; <_]6-�}�9ݤ��N���-����h�(w�7�y�zxU�~�'���o�yԴ�m��A���|^�<��Fџ��E�[�'T�W��U�-��W+,+��ˈ)�k�{�e�7�:î������6�Q[�$��{��@�J̆G{b��-ĵ���Ŀ�ߌx�t
�3�y�s3�g5�Ry��J��Pw�{=�p�th�WO*��H_�{����'����e�$��͏������M���h&zS��Kz����2���uU~{���`�N�ML.m�:|U�g?�A��������
l�/T�1�h*鵷�Րcfӑ����g'҂��N����5�����2w3��"�ThF�]�������T�;S��u�a�&����f=��V�,��)���rV���P}K{��~�`��E��#��9�O��:Έ;�Qe���l}wr|D募��=M��_W ���$�9���ad9��cs�#��8�����S0⯆\�\��ȋ�9]Ǟ�bj'�X�����w*�`w��Cd�Wu��PZ��畭����]�<j�n���)(0����_�'�̰T`{x���5S��v�L%�T�ۦ�</���̥mx���e�a���N�)���-lrm�$�^�H��T�-^�z%D���ǿ��w/��>V�{�t����L�w��BT�C�������/��SQ=!0P��d0_�~y��0u��p�M{E���5:Q��%:QCt���V��^�GQ�wV�{���,+���x���~�����{�k����ϵ�0��m5� ��D&Ja��=��Y�TT�Sx�Y��z�
~ω�9��t�!w��C�������,��������JJ�/��V*#�����-d����ǵ�ֶ*W��7�ҁ#�{��u��%2e^�q
�gW��'�5��Ƭ7�J����+������4��?�g��^Y� z����@M���3����6�`�)z5��9&����
��m�6��G�*�NO�󂤣E�M�K���;p:��Ԋ���[�e��q4�x����>ə\�Y��@��v��,�\H�<�e�!>���=���C=R�V�+��"�mzC���.�ّ�;ZS�V�o}�$m��pV��A8D� �9N'F�Oz�e
$��Hw�~�I1��'��v�H�J]V�|�C]����::J��q�V�����	4|��L�)��J��:M�0� ޟ%�=�nɚNJ��|�ְE��J�?>�*�LS1�M�.�y���(��E����C%�4;7�;B߭�&���:ۋ)�0Y�K��a��ގm�k���~�ݫ���?������a�����#qA�K¹,�[�\��� :�9���#��� ����M��̀�[͎��t�{��o�Î�R>Г����ҹ �R-���tK���R0�ߺ���w�YA9:Vs����5�Q�7mM�^&||zcTk6:�a��q�LO�4*�b��W�v�R�<]W=+̹K��M7('�!��Li��z��Y�2�`�T�t�/�t�̑�z��iV)��"����2;Y i�ÿG`�FI'PX��J�����=r�u4������&Ǯ�cBLL�
X�g�Y>L/=k��`:���'�'HN�����y%�ǫ�@�m_�8'm����e84m�Ͷ�/���V`m��I�<�]�l`W�+�e}��2p��Q9�N�=�����<0�w�Kϊ�����3\$	�R���/��)�BG��<^=`}�6? �Dz����+�ط���o����/P������3t;�XТ҇�W�[�k?��-�I'X����9��8s_�|��g��sݤ���t�a�]a���{����<�xF_p!�D���b� �5��?�ը3�����6>�H���?9��_�Vכ�ݧ�2/���qR~�?-5Ld�hh�=��k:�Q���#)m	��8�C�	��G![���h��(_\�Mk��ݧ��K��3X�?K:��~��,3+\�5�V�q�0P�J߈����d�ȴ�tO}�۩*����ܱ1����Y묐�D�j뷯]�!��8�*d<r8�>d��G��/���I�Lm �R/���w�Cע��7�.9�b��#�������:�X� ����������+_� )��9��A�)��l9�_�a;����*@iS���2����T`T����X���kR�q��Cic�e;��|� ��1_������)_��!4��è����)濽��9����:=7��s�1��a�y�	��9���n+�G�M���E�5��;��(����m�|��8�`i�5�Nk�*��4�
 _�M�	�>���[�a��t̍������ۉ��b|�0e��G"�\Z���a�R-���z�<+H0^@v�e0~�r|dT��q��˹�����aR�kࠤF������>�DpΔ� W��f'��"1�9$�q�ҲG�����3�����3d�SR���UQ���2��A�1dboS�X5���FbS���](�ȁ"�� +��.���ϳ�|���r��k�f��>�CF�+�ЭP"+����tq�Y�-_�*рY�5�?l,���)�h�c�U��ẏ�3��u�&��o=���B产��9�#'&�:l�M���u83�RQ�]V!���h=�4�վb��Y��V_�����^�=4Y/���j7�dK/�f8y�tB��D�#=�� � I��DC����u��O����������t4�j�(i�o��s�=��k��xJ�cj$�W�h�N/�xP6s@��z�q����^Ced�Zg�F�(U%�}``��2���a�[U��#F7�Z���=��ŚNb鞹;cQo��*8"�ޢ��V�(��t�ݙ�PN�VJ��d�y��%����Y�2����M���[��U���_=�����ѺCF�����u#H4C��������Rn���H��e�yGf���H`ml4�ƀ~a L�w��_�\w���D�K�/֤�֋�O��N��l����2��k�s�y?I.s�ek��?�ʾ�I"n��5��q"dn�u$h�z�i��o����w�rms���s]ANSD� ���a�������q��/[m�P����}����ZW?`z���WU���%X��~Ne�y�!I8�y�.�JƜbM��+��妌P��l�s��'*�[ُ��f��2��rM�uuS��׾	 r��s��
�)��PpA�|b���,�Q#]����M��\qC��g|?@?�����;g�l�W6�B�،�W����"}O�[��U���b�(CĜ�;_=�v��T���8�M�	B��2�ݰ�Y�_����K����8
-���m�_����.�奐��s8�G��E�1��z�υ�8#q�S١{c���ϗʝp�ҍ���p2o�I�f~�[�(�����`�%�e
)V3�<>(ǉa�l�	���SH�Xͱ�^��G������7�W�W"S����[!��#ް;p�H����L9�=�;����)!6M���3��suRL��^�r�&�F|!�@J|pEsx�؟�IB�h [�I^CBv��E{뷻z[��塅 �@Et�����w<:%6����'����"܌萸a�d%m��������Pc��B���P�n֨
���ʗ�f���Ǐ0tvf����N�Fϥ�俆�Z���Շn�p9�&���C�_��|�H?�A�]�Ob{٫5&,�����*.4P��s�0�*W!
qwG=�#Ry/������7�%K�����!��?�~U~�xp�#����*��齊uE\*&����Ё��C�ҭw�԰3J��g�����i(����bn�Zy#D?HӅ�|����D���om�.D��X&˚�mH��U�>X�=�+.Gw:��<K�8���)�w�U��W��5�J*���+'��8w	����S���6&��P�v������J�����S�Ĥy�eb��א"/�TV�.׾�9���Y~���E�}���ܖI�:۲4��<� n�8��MHպ�0]s���Q�Ϧ����v�|���E~������P(T~x���t�;�TBE�n�@�6o��Tv#6�ԥ�z�����QJ AH��.�C"�2�-��S\������\HR.��)�#���o�6�#{�`�e���c��=�����X3�@px�Pt@D�Ǎ�.�.b���soұ�*��@ݛ	�K�Ƹu�mA��������X��qt?Ӆ�Oށ@���/W�>�A�?�^�t� D�D���)=�Ó��T}kL$��ާQ&#�ZVs��Ѷ's��܉��Sw�MS֥g\-�?A�._��!ߑ���gP1��S��|�+�Ӗt l���M�$��/AA�ö�L�6�	1���Wm���U#x�ˀl�
�2;��@�C�S��)�.7����R��w��W��������@m?���&�o� z�F��B/j��k}:by�T, O�y�]W<�1��k��$j�s"F�'���sl=t�#a�޸����
����4�M�E�	�n=�`sQ\Z���tH�3n|g���[> DCP�l�
_QM����_�dB^��6��ɉ�z��aelv�"m�SCH��+M�N�K�np��T4��"�����O_����ASL����<H���#!�A��jTn��dP�!���4N����^��{M_�Lͫ�{����N7o�a�)��*z蛎	���`,>5x~��!�@�6���:�Z޾<v�I�[�
h7���,\*��N�yUۚkF�o��� �9�ٹL�u�o\���x���7�c�����P!�,�U���W�g�C}9�N�g��+׬L��FT/$𓈕L�@{��v7ӓ���v�[d�0�ǎ.�����:,bl��z
�X�0i9N�,�U�����@a��DX�@d��� p'c%~X�n[|�h#���Cl�{������A������jvZ��*��EW���԰</�[�3�=d������,Om�zA��j���E~Q?D�s|���dl:Ǧ�p�Na�k��P�������x!~@!\�����Q�}�����W�~?�!�����1 	z�R"=�3�$nZP�A�d�*�ѯ@��ۆT󭛖��h_�c,��o�(��|��r��r^Ώ7��0^�}���bO�1�B�b�	k4!0L�D#&����n���=��D�j�!='l�%�y�(F��2�=��U����5��{���N΋-ז:ˑ+�'��j�{#��(��0���	����E�g&���i���?p�gaT�DZ(�y������5��%��Q	v��z������x�������-P8�-r�pgU<o�h}�є-�r�,�VF�`n�R�^J:/�Ĵ��*q؈��m�٧�jj�bKΒ���O��I~!Eek�<J+R��*��|Z��/7��,�����"�('�tT�ʌ�����gA����OWq��=-}��\]�!�&�([���^G��
GM�/��־��3z��Zt��ȱ8q;�i�5T�����u=��A��O�O��]����ⱁ�e��������9�rL�����H��Ʀ��+1~I �n��CS�'Fg/Y~�s=�ػفZ�"����΅ḃP����X����&�8�_�K�ח[?&utej�Yގq ���W>-3K#P��dϦR��]���]�ժ5�J��a�a�����!#���!��q�S�F	fye���u��@F���-(J�0��+ܱ�\ԛO���XL��&������.@G,Y�u�[���94�<�C!\��h)�]p�s�	��u�4_��o�2�[��_�+�)1.�o�,S��5Z���D$c�=��}{�oȟ<���o1	���&�͍ն4�4���W$��x{a�v�[�OXڻa�"K�����[BCM�4(۠?�!����}M���/�/-�)�C?��� ���6���j`sh�G�-җJ�_�fo����z,'<�
��\�$�Hг�	'����mcx�bmtY�y��`�_���-qk�p���z/��O�"�!~�G8����.S���e�U�����Ĵ��L��ӿVC4�:uU%�+���#�^vf���]x�8#�ɥ4��m��?~⯘�ts���䯍aH|+���bV�98��
���?E5�����d4����_��ɜ�b�?�j
�e�B�;��,����:^�mL뚷��p�j-�C��6��B��`N�d��|������(.�H"PFmR|�ֶz�a{(D)_yG����{"C��k�mڛ<��l5�&�NKBΫ4���,c���WN4�����G#�\n�0�տ:�=�*mΥ�����?_���2�����ML��,�Q#1�jU��֐،�~�~z_�Սy����6�o�)�E��.�v<�h�zZ�����޸�YSn�>J+�}9���O��}}��w���ɀ?7�oS-rM}�#H��%JP6X;��&�:	=�δ*.I��`�i�d�2N�.bH;���c:[�1��k�v��`��⑲u9q��#h��V$%�o�i	�4�e#��m�;|\*`ٳ�e�e�a?Hc|Tý���%p=�/ ��Zp��'ް���΋�#c�=��8O)���{�	݅�ԗ�o�a�Jes%/fef����'�]�m���Ǯ���mY��s��6'!�a�$�I�oHd
�V2�O[K6��|���h����Sh�iş=Y'Ɩ�f�<�22�|�G-�����?Ά�f��%����!�*A��U�{V��ey~�vq�����GDG(�~Wo�9��F�����j� Y�?�v8�cK�L��7�L�6qoY�.�j��I���^�t
י�s���X�À��2�V=��B(`��v&|��r�1ϫ�n+�{]���
�r�b�u<U�>I̘��Ѧ�������l)�tD����ٗ��s��:`ߝ�JMaIPkcn������Oρ�E�R�dt0�c�S9��غ��9eA�P��c�҇�u��YB;NB��`�YOM�]�K�i����'�ϼ�^��I�b=B�������8�im��[��	�颂r����r{Ͻ��J�@��8ĸ������v�5�e58�۶Pa��t�G-R�x.R���*N��Ө�ǿM5�q�jѹ��,J���;WeGC,�gt��H�ǉ���Q�\�/�2p/�����[&�:?��(��ړ������n�%
���B��I+����K;�靺-��\Ƣ���y�v�s���Mr��������X7e����9*������rc��W����(����~�^�2��qqJ
4��o쓇v7�õ��E��j��D�2r����U���Ï_��I�?�B�jE e[��Y�+��#>6OZU�B	��
��a���d^�`�/�ۺ@���{}aL_����O�����_l��G�+���YO����λ�'u�dC�����)9i��i�u�7N��U�G���%p�?�~ׅ��Z����]I�(�y�PPC���)�%�mlm���u�ͣG���.�e1-����zd�\X�^��c����:��a뿞���@�+�p�x�����*w��Ԍ+l�e2�F4P2���@LJBAn0����T׎������N�=��h�R�h�_����s���QE;��S!��3�/��Ϫ��փJ{�s�|��Y=�:����^V˱ʦ-2��~�Ky��Q��Dlg���Uv%8`[��o�e=y�Wa~w�g4hɸ� �3��5�/�qT6a!��a��p����"z���W�OL��*"Y���w.J���^�Hv��%a��$d��ě��e �_'�!ߜzN"-}��T�{Y�D*Tx'H��\�3/&�)_���[��L�^\OtD:���.?����^�q�p�17���U�X�8arüOT�l���& �4��miR�����[�9C/��>�8��r0��ꇡӯTN���o5��C��ױ���T1.��*{l����6�ۤ�п�s�en�wK�m`t����d�o��Y�����ܟf���Os�j\ݫz@���~�7�w�BIE�Y�y?Ƕ��=�ION&�0EG���}�GG�M��e���;*A''`��ޭw���`����'л�D��2�0-�,���_ndO���f���;���4����嘆��gq ������P��9&�P��I7�̫ˤ�*�>\�|0cgV]����8`����^�4g�ٲ>���~������ER36�6�&G�d ofe�6���L�oR=m��L/��!B�N�K�۷��T�y��o�`�Bf��Ns���l���r;��,�$%w8��`��ڌR�����hl��������(O+�c�i#�F����������/<����V�{�_9r�K�70a�~�p���˧1mb��|�se�0jU?{�xo�Yc�7'�X�4	W�B�n��\\cDp�c^9IL��q���E��p`�!�����,�4W���*�`�w�Y��6["4��,ö�J]e�A�؟|� e�$�m�1�gۋ�r J;�s���9_�ߢ��_"W�@��wUp3o���Uk@Ė#�g+Rb�>+��-_����:a��_�Դ�!�* jmȚ��5I|!�ICT;0|���Dy�
�oV#���@7��q�b�5|4,t"9���Wv8��ĥgz�bY{�뽁����M bJ\�CV�����А�訤O������Ы�X�T�w���ȓNX����S��4���Br1ǒg6K.�N�O�����W��1�n��L���&BQ���RO�%=?��5
2[��g�ldh��b&}���f?v��{1��v�Zw��u�hs��bF27VO;ω4��X�G�]�KT���D�}.���/��0I����`'i:j��sC{�W�����c�%����+k+U�Ob&g4�Se���/��A�8�������QA�K��2�.	'�pjBrb拟�p�L�N��gp<��B���Zeyۄ�v��t���RO�Q}
F��+'Y�g�'��F���N��X��W�D68
�;J��9V�"?�?�"��Yw��p ��txh�4u��E���Ds�����K����V���(� ��XϏ��ݪ��Y\��f�bï���'
��ܷ���B⪣�$Y]�]���0jf�z�d.�%:c��Q���.�>T�-L����,}��� N���.�bn�7���]'���v��7���ީ'���Â �*����bR���}����#����R�UG�,��b�1��#��N� `-��}i�t�u<�ܲ�.��0$Q�����y6���C׿����g�ge�XC�	�4�c�E�����&_-��-�D���5W�F�1��w�;"�ۢ�𡎤Q\7����йd��_HSk�|�_��U7g�!�[d*.7m��&��;p�.P
��r?6a�/�A;��R��l�S�A��-�tD�p�U*f��C��wY`�>�fN�H̰Rll�~�o�'��3ko��O͛c�w;��"�������x�Ɔ�D ���1u�����տ�(C����'ۅZ58���Ż��k�u���-𡒻��bt@�����'2��B��FF��������R����x,f��_;��z'O���W�!�汎��K�:����7��(�}�&�ŭ����wsx`����iDP�[ 슺��/c��Z�e����y��a�D�>���z�o5se<�o֊�'����-�������Y�)�p������߮�8�Gg�pe$ݛ��^[�[�Mw���|���>_�޹��'��[�]M��/~��G���d�"M�4��5Or��OV(���=[�D�0_Y���m�~�`����*�T��1�lX�.0�prX(<�^�������Htu�=	�v�uRY��E�0
'�G�5��?O0}��[��jJ�5"&�P~�F:J�G.a�?l,�����jk�A�� Ir;�s&y�й�ɾ���_ù[��t9�:�w"=�}/��RăT®�"��_���g5»���-xᯁ�1�h��O]��EBy�<�X�
L;�{:�4Z�H�n{���E�F�GBM4LvA����y0ܩ���d�C�T�贐/�bYē���L�	nu�5�Mپ��%@�M%F.����׾tl��r��S�j�0��+��~8�$em�y!w͕��`*���%�&=�����A�B����؛��jU(����ׇ��T���]ӿ8�3��;�pz�ss��OP6�O[�2����tLz�J;�?7 ����io����[{�O@������m��wS��~}ie!�/O|�1���gu�� �,X��\\�IŒg�O9F4;�ǿ�d�@J���SPބ��W�zx1L�m�7��Ɛ4�;>�b�J�=s�̿���ҝ&��eP�q�o|R�K�*)a���nC�����wY�����T;N4gj�a%>�sLh�t�=5���)M5��|��B8��f���h,2e��k�O��+�l
��Y����Ox��fmŦ���x�W��'bS+��J)s�#~�`��}ԃN2"�Ǜ�ő�E�d&�kH�x)U�nL���Y����Or3���C�/�,��Z���T!`�~�P��R+P�oM�����¢Uw��E�3R��U�)~�<1���Ga/���9\��weQ&�~�����E�k;�X��Xn\�).��J>^��X	?�LXM�� t��iӘO�œ�����{Y (���n��CӘ���w	��RE��c���c���s�o\�D�4�m���w�!���&���Ӛ'�M�L��UU俻�@�����_�a�F�#��ӫמ�Ŷ�πՋ,�!��4t,e�q_@s�M�4 ��+)}/�	�u�9�!��̾���A(:JR_�;�۫���=0 ��"}SJ���Qc�6�BJIs��+��� �S�«�^{��B�=z=�uq��l��<ŠA}_0�%���Ì�;�)��z.I8yǌTlZL�,'��ȁ,�3G��ע¸vj��<�I�����v�y����sB%բ:1e�@�@Q���g�'�U6Dh	E�Ov�A��1�O-Ͻ�兺$��c#�.��c!M��'��K���ʸc�+&����zK�j�I	X�6@gR=<���_��h}����^��X��hw�"pN�i��:}����qhڀ++�;BP4���i^��*�}n=�O��1鲡K�Ew��GG�h��6@�f�i�:�]�s�^�\�RJ�4�²s�5�E�A�f].EWen�3�#������8]R�R�9��KT�:��PZ�`1�h����wO���B��-U�(��l�Y��6�֥u�S�	?��y��_��n��{e=j�4�fc,�Y<;-�8�,�[�'����d#2ׂ���=�/�e�v<�o��X��8���)��W6j�O��s:�P�lg2���%���b���מk��x�|��Q�A��Mz��m~R}-���)ب��{��揝/`�%�׈8�ܣ_�8����<L|��W?Kp����*#b���Mc�y䒆 -p�� 5��`��uoK��T��034dHZAs�p �
J)���'�����O.Ȟ��MV�%��9F#_��J�r��{Q��Q���w�^XZmh��֚�ߑ�\��������6.���	�c�1G/�����=[�e�p���Ad�Q���{E��R���h�й��3�&��j��d1�`U��'-���G��z� -��C�/[����5�m�{�r{���ϕ�Ir�\C`z,�x��,�$W|�;)z~C	W��v�{_�ycx�>�D�_)����=86����,�;�xFAp6{W��F���]q��ࢱGYid��A�,E"ˇ^,�-�)�w �7ɏ�k���$�B�'���Bs�#3��Y�_҉���:�f-yv�`�����$�Na�*�:g��r��pN��������Y֤����b�L�h�P}-�����y�c�aRe�?��Wo�[]����ZS�����0g=ʁ6G�PK�K F�=%v3�,��HKCŊ�O�y�|2Ԡ7� ��8��>K*^L�+Q�����ʵ��'}�J�|cQ18��<n��bښ�
�{8L��|���|[��މ��p�֙V#y�5���&ACҮ�!��_�ŋ�	W��yVd�4{�u�aD�Lh�T��:��96Q��Ю��'� Նl(�V7�%�n��-�Vz�#�zX5@A�������ӦV���p	�!J��d����	%2^v�}mlQ���Nl8(�(��� @�Nd���;W1��k���O͟/����u��t�B��s�g��1u$a-�����o��v�0�8ZZn�I�ȪL ��}��+Z��d�ϗ�5��H<�yc��yiY�����5{&�{ޭ^�nD�]6[���W�q"Q9v���ٿ&���G�_P���"�ڎ��E���h���}mk�b���TYQ�#V�[�ƀ��W�O���_x���v�BK"�-#�>@�x�W���;�%;�@B�1B?a��)���_�������s �9��ƌ���9�Y^�������K��z�4����h:���B�?�%͕�ȁ�,{63��H�D2VK�	���1�td>�ybAz��'����x99��N"vjP=T��?�H��[Z�Hg!g��L�Q61=�������b^��.�	<nk���XRZW2n�$E����LW�ӫl~H�crJ���WQ��x[���Tel�j��	���9S*�����*Zz	R��8�/�pl�����%%�W�֜���\�F锂Q�q���2�d�k�4v+)h�����y� m���Nk�����&) NE�ӎ�����S�X�x��BȻ?�]Ε?7;q�3�<�gIm-� F&-�(��ݫǽ��$�@�?X��,���s�$�kt��j������d��_FD�R>_*絊����Z�޾-���2U�h�dN�Ҁ?z%��K����ٵͪ��Rj v�l�9�ߵ5;���p�1�����o�`K>5����g-�H�ITrLQa�9�I������o_�wϗ�<�mX�	zx<uIO�XÝ�����I&����1Ԙ�k�G�%
x�t�V�R�z�x�����N�~2�� �g�߮ʻY�Z��CǾ��j}�����6j/�ʊƭv&`�it��q蝜BT�s�<?�w�x�b�{��7�> ���}�Mw�6����0r�W��h���g�[5>%�*Z�EKd�kF��7P~��5.J|:�F�x��$����>�|�]Aw�w:�d���Ŀ�����F��<S��sL��W��n<�f�(��/ߋ�g�pP)v���i^�Y.K ���i��g�!u�UD;��/�ұ� �g�
$=�㇈[a��B��VX���S�x�y����m{�H+t<d��~� `�G)j����d�U�@������wp�F5n��pW����s���o������h|j�:�of��$��t|�<~���Az�5�k�vcWU�q_Ѡ��l^8��kg#�n3�5�к���2s�_�����r;7�!֨�uPO���'RQ=�����������i�m��$���ڍ����v���=�����u����M���#���v�agd����45P]FCp��3?�\�&?�p�-�+o����r��s��7�{��pPn���Zc���g�V.��/ǜ�#3��(�N���}h\��[����3>��x'���f����LHX��k�:2<p���%c�c�TO8����|	�ahA1�V�� ؼK]���v1�ی�X���~}���k�x|+�E)(��G}N�H��75�T�n:d�눕�h �n�D�G�V�gmc��!4�v3�>�l���"�>nB��v:I��$����>����Bi\���.������]1k�F�V���ѺT�zB��tY�P�>b�������:9����}*b ��;iY�9�1wwm��QrƮi�c�5?�Vl/��I�0��E�[#���-=^������_y��x���
 +M�J�-	�
���'X�e���3�?/�z��`�
G޿Tg4��=��үO	��db
�Ek�K�C���8�������黭����n*����Ĺ?ƿ�6TF.?�P�4}{�K��yhJ�{,o�E%���r;�wO�Y�hl�v�$r^	ډ��Ɉ�y �.�
�#��2��̚�\��҈��'��7��vV���0��ڤ�����* K¹b�+�w��7�][q\'g�)�A��ޫ�)��T$�=b� �۔.��q4QU�3�0X�p�E�P<s����&圹`����� Du�Lv�M5�)�V���=n�q:>i�gW��ՅU(���Bf���~̭i��%)Q��;�@)�B���|��k���O�Fɻ`�I��V�S�Fo�������y�G��!��L�C�5���o����G~�r?,8��K!tTG�G�8���Z��(��̖=�|x�lG��y�#�R]Bv�G��WFb/a!�yQ?�V*�����n��95�A �GS��j��w�3��r�viü���߈^��g��#$τ�Z�י$�٭� G[-��:a�r��3�����&�W�@���Γ?����qS���k�>�������֣th�����D=�%�ɢ@p���֥L�У��R_��q����E&�o@n��BOԏ����'�?"I�`&쇪�_������\�v1�H[Ӵ�8	ƜGPWh�K��`+P�\
g���Vx���~"�lܦ-P��ݺv���LB��@��~�$*���)F��	=��#�rb-�1Ѧ�
?Ͳ�^k�����u�7��XG="	�;z�DЛ�
pq�h�f����V����_�}��ߊ;Gǭ/8J%�!8�-^��A*��~�Z٧+��|Գ��gԒQ�ł6I2�Ж�$ž��4Nd�����I��������sܔP�k����<_1�`(�U�7���@8�Xߛ���V��8���e������o���Ï�oi���_D�i?1*t�KYk�W�v?���� ��>���,�ԣ�B�uݪ��s�2�o����S�,������6ŷ�e����*�97�D���g���֪��i��xT�T���c;�!ז�_	�MB�@�	�_Й�$����Q}��JH�ۖІ2ⓥ��K�c�;m�)csO�Y�u���;�2��>��2��N?�B��ZeQ�<ǭ�r K��U|����6��v����Ye��ſ�p ��9C;�R�k�����n��EI�]h�b�pb����?�16�����l�����P�ۛ^p ~"�HU��z�r��K�w����l<�ol��6Uy�X�SSj��)5t1/��I��.�N�S�.���3���/㼩�?�~���L�l<!_k�x�F���k�ppI�9iQ,�)N�v��˾�٪$7��9�);������NHJbs��cp;?��g~,)����F�j�mG�<\�2fv����+�*�v��c� ������'�n�j���l|�d�T�G3�ҧ#}VI�$��&�K�l׋F i(n��\lh�  0�\L�JQ\KD���w�U�>�yNNN�O��k��`�~�����Х��Vƕ2��6t�Q�N�~�l���gCw|$	�NO�:�'i	8�u��A^��Gѽ���DL�.�w$ *�4sw1>/�r�-�L��G��>:���:o��~���@-h�뚸^[92�a蟭E���m�C����U�`�fHj�7t�Pd�)��@�<Yw�Q7��	 �'B�>�Qv�9�ʷQ�7�<д{�U�z��/(2��ʼ��?0$?E�7�Vcm��|V���ۃ�"j���0��	a�\ E�|��1IK�r���d����h���j�m� �f ;OY��Sf@Q��vj�H߷��a ��(f�Z�g]��}+&���N��%!Z��t��`-���2N��t��#�f��_=�fq�̣��zrώs����|M�n �L46ن�L�t����T���Ye�&����ʀ`i����{�!e<D�&�^6�.�]�"���� z`蹅eÂ�r�z��ѵ�E���A߆k�j����kp���X����c������d���2��{��0���@'�q�M���/g�L�2>P�g���<zK�%��춋��($
��Cf^�X��<ۣ���u��G��cZ�MZ�[Ϗ�z��h ~^�z;1�Y���F���{U���x��*̯_T����|j�_0�D5��;b�>'�h�,s��������p���w�����+�i�[7!����|廛!�]�j�ޒ�s�����ͷ���̟4P�^}(�ܴT�7ݬ��!A�I��,����N) �k���%f�A�G9^�zT�ҁy~������u����:���>�k�1�0֠���1���yv�JTC���IeDS��xVo�f-Z����BX�����2�����'iF���s��|ѧ5?r.�2~�/Ap�1�~��=H'�u`�ze&���U�r��C},�����IV6�y�M��f)���w�fDY���2���EF�����wE�v�Q��Ժ��k�����9����*G؉�b$G+U�yρY �(;�D��D8� ��G��O֎�����X>����k��7Z�kFj�hcӅ����S�>,R�d������2��m߷�ye�ks�zk�;��c���E��T,Fx�.�?.��9�:�=������ad����u���9C@[�B�g�ސ���*�������J���@��9���5X+���.D�v���)��g^����e��������W©�'����O[38�5�hK��ZCr�1�����3�40�B$�6�a������#�% �\��\��eM�yk��a�ge�w
8u\A1ډ>�sV.��V�g�)���=.�9��.�/'�B��)� )(�J��\�/9ߵ���*�7�B��!��w���ĝ���J~���0 �l�5�Rc��F�@�M���V9/�a�ٲ��U�)�����=�~^��Ë��X��aC|�����N'g�� ��ؗHmuWݞuYd���ϞFy���^�$���{�vݯϖ��#���zP������������@���F&���))Ο�u��+��]��!G�cwE��
/9k*$�[k+�E�j�u57��_�s�Q� �(��ׄʓ������p��������o�/coF��JJ
�E�
�S�>��оߝnr/�>!!�L�1����t�>�\A��@֚� i�L�3�b������Vq15�P�}��,oF}|�fǔ4Qw��#��k����bnZ[���L}4Ҍ*�a�B~���V���Do�\��OqeƔ��Ӽ����|��ײZ|}��J�Ƨ�(����7���s���7�ᘭU6��i�!�v48���׻�O���uh�´�A��3�64�F��A��C�	���N��o|�����^�k����9�Z��x1�OQ�[�.�Xk(A����,e��]֌F'�[�ÝbS/�#�?��*��}D�"eЈ��H�tyQ@�;�E:�NE��.�J��E������ ����׺��������}���=�#DX~L6�Ng�eY�K���B�j ϯ�6����I/�\2~�|�cp�j�/�ܝ����-z�vIm&#�{7��sWR��82��IFq�,���\�ZJ��Ӷn� u�q�w!����!�)îO�M���JJ�8Bx��H�aC\�Q5��%U�$�Ga���<�[XIg��J!t���y�<�pzvT[,�^���4�T���z��j�$���d����!H���R�9��N,t5�o�c���3�����KɳMd16��P�p����>7�����lӛ�N�<�28���H���N'��_�Q-�?2��u�f�y�x�9�\�iB��У-//հ���|����/Oy�t�4ڗ��Bfre������0�l��}$�\2-gh|�%��荆	�0-���j'}~{�b|{.?�a�	_q�ϢH��1:k��t��̎��^��]"x�[Y�S��E���D��U�Cl�wm��u�U#.5�_H�ܽ�oU��i�)yI���(W��lƦU��Ky��0�.n��$�D��c��ݑ�5��D��9���)JVI�6�Y/g��Q;�g�l���-����W���խjww}������-��$x�϶a!�ې�>h���ߊF�a��TdM����}�Օ6n�>4졸����ȼ��9�8�j����^��7�S03���]��U���ͮU$���`c�<`�?~z��r㻘��6��XW�{i��V�|O�Ӓ�'ۿh� �*�[�L��=.�D��@�w�R�#��VJ����������ӿS�]�N1��E+&�f��͂��N�i�ٖ��m�8��%��E�Ců������_����؛-�v���YB�vZ}q���/rQ��>����q�@ާG��c
�S*ٛ����%�g�I����kn����Ţ4�$*�_��J����G�[6�F_�d���WٷwQ�W::Of��p�9��.���/s���gou�WEh�--����d�C��j������6p3$	�C1T	�u~)�k��\i�˳&�g���t�b�h	/)N��1pu�@r���F���0y���BC�����?��,�/U��ZZ��(KW��b�O�g�6I�:CƷ���{��1�aʑ+Z���]4���>D.�_����gD�谏�/�l0�'�x����G�A�#�xg7�{
�O�[Y{���M��[����#P"$ـ������a���o�uT5��vS���,68U��6��m��Ƞ{0�Yrj43 �]��,�^��rA��p#�k�;�����Kg�	¬pD\W�Gw@Ȯ��+Yk����0��.G�"�s���~���=�?�`�	R��k�
#�:DEv�(��G�~��/ə�ND��.��(4�ӓ[��U�m،��P@����j=<��ks��R��h@�VO����i�HDE�T-��;v����r��c�J�U�/�9��	+i=+ M���bYsv���k�zT�!�뙈vz�6��5ѭ��v��]_[4���W�jz�t!�G��T��k� Lۑ
��I���d ����zK@���g�LD4��n��
�6}�3��}�['"��v5j��Ug��_B�ڹ���D1�3u{.͓�^j+T-�/]�RV�Zd�웟�V�����c�L�c_�6s��ׯ�"۸�Hz��uU@����K�]������j�.�P]�'�V��N7�ga�<�O��ӒK�X�/3lg��5�±���*�cd��BVul�5�d�l
=�K�f�mzyr���L�
���ZZ��h�Rj.��nl8���҅g�+��.�ޝ����u[��.�gu�g�x�S�6]���ߩl���� �n�l�o�~="T���ùR�'��?�rú݄�Δ�o��!pm�'�����,���� 8�q�l���Qa���յ[�nȱރ�X��t)S�-�nbk7yKF�*�s=P��Q��z��4�h�����`��|����pd��(ӲD'��߯�m����D�x�����@����&>����P<��,�1F���3}�����Л"����#X�������'���JG�j̜я�K>^� \-\�=,������b��.8���3'�mt��8�{�ޘ.-'���uWƍJ�ˆĥV��md��@"k���h�u1��K��Ef������V��v�p�f|lRn x��5<�QW*��K'�@�@�ՙ���j��	1F:%�C9����wPt��{���R�,yW� ���͝w`d�<)w�LÊ���k�9�օ���ԩ�U����U�z(A�q4:X��1u?7	$����	r$�0�^��!��t�S'�)}���e�WZt�����O�5�CO.ѧD^U�KJ˯a���j���8c���cQ��u=��p@���J��w��S禊a����n��w�5�bu�]N6��ҁvs�Z�f�yt��`��X��:����vU���+6�|6CE�O�կ�v�y�Աn�5�g��S״L=h�Y�%5��c5�g�+0�߈�"f]vFz��V���̝:�4��6�^*���	��&�}Z��8o�����v!�f���S����^�'��؋�(��uB�����,݌WF�"�J� %L���Iv�h�v���Q���08�h�T��%^N������VW���"���9�2X�s|����f~:��+��e��/.(���Lɛ�Q��`N�x%�v,_�7qf~�����Cl��'���2l����I��)�+���ԩ"�D>$�h�i؝�]ĭ���t&M}²o�*v�Q^��\����׀����j
�>-PCp�<��������q������H�O:��l��x�X0]��y��a���m��=XH[��<�jtqW-]&EF���g��ATp�,/�݀n���3-Z���;��n4kZ�TP.�(��]����?��A��4k���Fk�o�<�"�3HC1�F� �a鄙��Q�(��[���}��,�5�	����Q����4��g��ͤ[yӑ�@�k;]�.��-�t?7��J��Zf�N>�jF)ƴ��}���~��<����Q���֬	"'��mѝ彩����²�P%�ən�G�,h��K����@"3���Mlq��i|,�/l�anj��@����E���VY�uW��:�J�̡4�S�S?�P���%��l[�g�k������ڴn�z%����/��N���o<��ɪ�[
��J�+ 8� ���-�Bm���QKwoծ��du����$���F������%�� `\�]�XkN	�ߩ$ ���G��}%޹�
凷S�}�Y����O?:ڵ�9V���N���X�>Md���f��2����s��hx�����E;���=�Oċ��^�^�g_���w-���H�g������uy�a"�K�t���BF2���Ҟs"S�p3^�\�ǁ��6$&'V2}�5��\�I&�+�YȊ\�E�]�:�d"���%m���>W��t�@�R�j�>Y^Ȏ��Jli�fw��K��=jS��K���;�Ư:쌑x���#^G_�8�Dt��3��#G�@D��>	�%1*�+�U?B_,�^.R�NvxгH����?%�r�{�I����3o=e�l�48ݵ����ۢ7��oĬ���aO��N%*���(z�R���Dm<d�4M)z��ۧ^�K�)7W�J��>f��c���kX���o�lRx߸/JV��g��Y���Z}�E��=a��-��:)�V
ɾ؏�j8��朒�l.���5����d�> �f�/]�o����q���&�|k�!�W�<�����ʷb�l8�P��u��W����
��1n|�J�韨���S�݆�`ś���>��u�}6�թ�xN��`��q6����w�|Z�%/��C�mۓ�W�?v�U=��鉜r�A~�Ø
��Z�bU@��ji���}I�`��6�q�/�0if�MlX�]��??���Q�6��<�h"��k�W�5\�b�o���-M�6��A[��׾�w�����*�Te���D����2+_NKw��VVzIQ�;-���
��9T�&aSi��K�rZlM��c ��XN���XF��e�Y����Rbb�����O����f�U]�)�)��:�'���T39ߑ+-O�v]��IB��2��u�h��.!����G�&�����q
լ#Ў��i��j�u��"�Զ��o�1qI��S�s]vX��4�g}�����q��K	���S�t�5�����������"U�L��ri��/�<�raq�{Y5f�d&�i� F���OL��Z5�-��
�7��VZ��нJ�V͇�	%*Zwqn���H'������	O�:g/7�d ��N�ݲ�����6{~���̫���8c�"Y\^O���]8������F_���g����E����^n��2nT̔��������j�I-+1K^�1���홿\O���RO���W��^��y��I��?$�3<���KΙY�n�ꗧl#B�XM�pKhUG��^�t�Q�����h�t���˕���n��as�-��#�`���i�C�ua`(�p
���C(�Ȱ�5�%n\x+  ��O�#gj\�Ej���K�Ԓ+	��M堥�~�`��e}�V��U�j�����䰿�y���OjT+���Eڱ3*p�/�tdӉc��$r)(��6 ގ@�4T_}ڽ�'��jў&��7�D��?ۦ]�j�m��%իh�-V%�������}�¿|D:ǟrgNƦ���z;��3��E"Ζ�q�/����0:К���TN�6�3���������>�u���!�{��F�L��n���`�� ����U����v-�5r� l46r�ؘK;z�b]4�*!�r``�(�1գ�i܄_n�U��U�i�}�0�4��/���r��I���ԗ���G|�h{�+=�M�b���E�*�Q4�y�{Ұvݪ���f�	���0ϵs0Zya���tu�q���&��qIC���T�($.������H��3N�_킊�*�v�g����Gu��\3�����Wx���J`���Τ��Q�֗+B���.wY��6���0�v�Y��S{�� (M%��n��Y��+���`�E=�$��e��Eö���Y��e����q�5�YUo��?��Y�l��8\�+�C��x�:2�}א���(�Z�?~Z�}ja�Y>��ϏJ��y�f�����5N�n��^��@$�_�	���:�T3P�(ċ𺫰}O��wk�����ᩩ��t��`Qgcfу@f��rm�bn}T�/�4%8��o��7�5�t-۹_}�JD��������O�M����v����]��u�V����w�(f=|9�|Fn��s�(��$�T���!�g}��+Q�^"�xܷo���k�m�%\�T�M��� ��8I��W�&��}U>E����+Fw�,�����5��';�@:�:q�m����Ł	��/�.�讕�Y4�(f-�1q��ƫ�}.�n��v�J���+�S��t��~$�!����Ŕ7-�qAF\��i����;vk]�8�879�V�/��.��q���zx�j�f���q�y�j�ԣ�t�G��3K����M�t��n�'P=Bf�A�[�}�Xm��(d���O�R�����S��P�	{H��(��x�����C�=1ګY�G$��fW��ɧ���!�$��w��FڅQ%��o�x��\���e�vp�>�r��s>TS�B���Q�3��I5�^7,TRL�|{u��m0�1�l{y��Z�y��?��dĬU���Ԯ>/u:�ɒ̔��^�j� �ퟌl��p1�^
x�ޝ����i�8.�=О���O���{5������0�ʼ��KALOEBOMq�""���*�b�,ed�m����G|o����j)slW�Nh���L��Oy������\���~��w��r��~M2SsU��;j���^K;�XZ������u�"����ޚ=�e��U��}�8�.���+;J���X�� \�^����[��kF���b���KB�k��q0�6�P}۵Y5�5��l�6��▱t-�eG��5�l���ژ}�\����}LҬ��V�E9&��m?)>}�(��Uƣ�;��b�'���gW�:�qՓn��/��!l\ܣ�3
�Y�����[���+x�Ys��;q�\g�Q��"��}��)Ib�Iqa��&Ȁ;�����H?��{C�Ϟ���Τ[�j��6-w�����V(����u>��� pE��ܞ���\ }���68s�p��8!��m1f�m��:[d�0�p��}ei��=m֩5�4?���v`6<:��j�^ߙ��	q���6�g��!a�@�p	{�O�Q|8�#*���	�U�����z�6h$�1�z��mC���������E��>�7����9�����G�Al���?m��G`��S���Ye௵Ƒ�Ы�m>�:�31Ia2�߳��w.?���ڥ�r��k�qqU_����{B|���(����j�8�K��1u�~o��o�W��3�w�	}f \iL��l� P�y���x7t�(�X�s�J�=j3��
�S�-ksg޷�4�A��p��-�0�ʎ*O( ���K�R��Y۝��j�F���3�dk&�Zt��t�ӣ������j%J0e�v��w���������U��s@��Y�z�6*@��=�z �ѳx� '$����z�k9-����M�TcA��52��h�"1�9y��6X�jQ��SG�"�E�!�_@��^C��u�_D+$bjͥv��^��M��i�1-�i���5
Yq�#�(�V�䁈�P��l���\�gVc�u��S9�%3hMf��
;d�d�UG�SM��x��<��1��Y)�eĬ0���G����S�5��[Ѓ�i��l���h��3���Q:�]�Q
>r��&shn�b���	Ki�"s�]�rx������[�0&�qxG���_���5�z8`�w�3`cU��g�ɫ���[�	2�X:k�.(c��s�ܔ��-�p��h��* ��+ҡaV�Xº��Q|�ފ���fr�eN1Fw%#~o�[����_��R�[�5�㆝�>�@�(pcd�G�(�3t�H�m���#@�u\����=���D�|D���dݪ�"#fl�b!��]_U���a!�Ƣ1Y^��a�)!��c+��:��p�c{mKne$\�B쳸��5���-b��mxJ
6��l县�*�A���|-R���Cycږ	�n�G9fC�s i}���#�$z��}�ad��c;R��QCr3.fq]�6tm�U;>��rt;�;�"�G@�?�,п���@�w!���c�X,e?���򉨛T�f�jN��T>�����V����?Ct�*.ʬ+k�����aU 8<Aِ?���İ�W�]�wl��5�����5� `��*̲�a#�s��<4o�x�s�d�Ѐ�엎�����M�}�`L��9Q�~ܕ��ePA7��*R��g��& �.�!G���?����]=������S˂7a�A��!�?�!�� "2:�De���C����J��P������{9~��ʣ�<ގ�@'�?Z3�Ya���X�ݶ���ڟքH��(m�&S���9���l�fLH,],��P�?����n�$WJ�ʑC��O��ח��;�<�A~~t@�Г��q�w�?N�
*�T���]��M�P�3Ф��E�E�_0�[���؁�=�������Æ��J6���)�%8Rt��:ݫȑ���|=���R��߽��x��ޟ�ͳQ]>���#�|�CnZ���H�c���aoy�6'�L���t<���!�F���T��.�aň�}�m3��v�t����}菺��ށK�Vo������hZj�\������|��a����� ��D�4iaE�v�f�ĘD�����+�!�Y��: �V(�kb�4�����XA�b��_��L�K'ܐZ�wF�����H�ʿ�*�r�4�hl��M�_yÿ���v�g��SZ���e%;MNe !��A�x�q�:�4���׌\���[e�&�@��I�4�VC�lK��a=3�.�7�E�N&.�E**|ˑ��`[���o��T�\��s���;o�Z-0�(���&s�\�H�ge$�+�f��@@�$&��g��U5�f�A��e�1���;1�6ĿO�� �ޡ�+����ˋ�XX�Yl���u��:�E"q���0�R�-����m�b�ӫ��}l�!�����g�ܚj*T��HUz�N ���~������Փ�ak5:x���y�I�ߠ@i�Af�.6r>}�w��l,���'�h��}c8��K��ܵ����i���]�oq�3+/Md�$��}�[||��,��.���u�S}�b�Ȫ���g� Z>����m�;������z���n)�w��V�]��t^Wut�O9Qs����N��s����C`�=����CD�����Y�#��Fk�Q>#8���������N&���S�J�/<��fr�g�?��l'�c������m�$���_�sٳ|����8����f4�ʼ���V��G����W����5���;B��{2�L�t���������e��\*�2Z� ֔M�"�)Y�?����$jv�F6����3�Z�p5'��}V�'��*�(dd��� �+y�JG��E�:���;DR[�%�@��n@��kc�����r����A.��1XZ�d;��f��O�^6��xM<��D����xlG�e5h��R�E����*�A�h�'}צ�`z�-�%��H�m�*��u�(W�v�ddzC%�wq�9*���V"�̭N�c�}��*�gxU�.<z.��^>g��	J(5Ѽ�ǉ��H�YNY�Y�XT��h���D���"�k�+��8� ����F="�ڋ�1t|q�Y����a,�5㸟E+�u>�3r=A;���"���l����|	Ød�ёƫ'�_����d5�F��g�<J��+ϗ�`r�?؟ECB#�u]k�d�,lbpt�k�އl��첄�ʘ���p�Lz�[�~ؼ�p�?�w'GLϊ�]��e�b��+�\1K"�^�:B&���{�>� �PRS�2�0��**����<v&YG{Sŭ,��cr�P.5�qW�E�c2(z P����NuGܗE��@<�3�4K�߱��1������߹)Y_���[�c��V��RY��̞9[�Y��H��m��X�¾���=�mV�gs:��cԛ��5�����'�iÔ����(WNz�����]!�s����6�{r��ߙ����d �,#������
7��#��;*u�z�GC��HE�U5�8+�awf�`�y��i*��nT��ǡ�~��O�����E��>��V �'��6�L���Å����W��0����xZE(#jd��lf�פ���M{�����P��>n�#-��X+V���Y����1�����(|����?��o����L�'ƨ�b���"��II}6y���EM	��&�k��_	7���"� �l7{P4gA��xw{{5?���&�]�^�#��nG���G�͠q����3*puxݳj�H�<�7���O��12Z4� ���i�Kzt�6�
_6N�h�z���9t#Ȫ*�� �
f�Pڭ
�PZ;�E��
)��l�!|B}@U�F]�w��J;��c������{��aBj��$�(�2�V]����{�FW�l�G����ʧ	��a+߳?h����+��g_��<�����7���GO��.��f �H�þ:]d��1��x�gc��5�R�Y�^�v4L��O�,�l�д8隗3�E|_'m\���[�7n�}Y�u"�J<;60�B9y��jß��v�A}L`�Й�E+��_ڶ �]g�H�����Na���������s�WR%1�A͎�h#��x ��V.Z"^"�X��v�*�a��P��S��S�9�> i�۔����>"U>����ᓣ���=_EW��Q����פ��,�sC@�O=�]������:�X%�f@�V�7���.<���'PU���)uIJ���ŭ)V���g�`V���	�d[��ˎ��"��O���&�r�6.��E�dP �s��h��ֲ�:������h`&�Aѯp�yd|&C9T�w�M ]~�c97\����g�n58�������)�z��w���B�қ*<?�yn�&
�]�wQ�#�ƴ�i&��u��^�ezѵ�5?�V��u3ࣶ����޶O�.�a��g-꼅����:Ì�߻�Ρ�ye$9�ށ�> ;j���`S�4��s�w74ˈ��"+7�(�ny1z)�	7�h�d���S�7f��|��z�k��l4���? 2:�?�&��4N���ox^�N?�ͤ�q�8cd,+fD\��;'vA+y�Ť��/N�{k�p:@G�ס- ��t�U+����]�y����x8��Ø.����`�|]�J�Y�~gNR@iW�J�Sv]GeĈܙAܨ0{��i���f��y|Є�@�ޑĤ��T�1e�E�6�U�T���H?~�ȴ�r@P�(��>*0����o��y��〼��m�r���A|���@�eu��kY��`4_����D>�aJ0�}wc�!�����q�I*@�Zz�mꏠ�`��4������$����N�rS�H��޺n�o�O�ܿ�.f����,�������@�l�K�5y��}��~�* WЄ2�~�~6��I� �������Z
P2G��(Q��7>���J�PA�����OGn�*�������Xej�������Mp[�>h�[�L�E�-�_���f[�S�
��E���?��)�7{B�6��0U�n ��;X�2�5N�<�M馓W7$��  �NC���B)��b����k����7]1���X0�߉%�`���ߓ����D��1`�r
�4�:W��?�w����G\��{o�~ ���F%Y?��H�<{�ccW@�� �W���8,:����$/�p5p����le̦zx_g��{x3����CV`� Z�πx'����f@�BZ���_�c�B���݉4f�[����@�����,��O�>"�����?P r��{����/���-�w�<���9���AAq�	�Y�[���sO8��M�!W�~� ���c|t���xFm��LɊ�2����{n(�Pޣ�<�Q�H2
�H��}���y����jϞ|��u��s��WD�{�*�C�Y�D�B����X�<���tS]���ׯ���s��M�����O��y������Gm�l-�Q1H�e�_���K�TB��E\��D*%�Z�l}�w�"���8���ȯ�Ro opt�y�箣?�{{T���E��,�r��-T|��Ro��1�is�V�yK59���n�n���B�r�Y��? ��.i1Hj�'�]��g�f/p)�PT^|���:��wlF�Km�w��w�$�b��P�9�ȕը�AXo婎E���C�@G����=�D���T���w��/!�T,����ӕ2a�L�w�����I�;i�P)Uݽ�{��(�|��̷yRP���"~�с�`��2�%/����Z�XVD³[|;�� Es+���)? �Z/C��q�'oo��X-�a�4 �n��I��`�	����BXP>#؈�9rZ�R+���w-I��D�^p!]���#��J ' '�ga7��܈��'<Ac���|�͑�UF��-��w�b��4��.v,�Z.�X���0z�g +n��g�3~;G�I�v�^!��F�2�$�.f��0�*I����"f:�:xU�'T�8@3J ڤT!���J�P�v=P���������	u��p�\F������i�:�A>�ug=a��]z�V��?7���Ř���BxR��g�YInA��I��a��)rL����s�]�Vh�$�t% nD�w#�;(��a�������t�$%��T|�խ��Wjl-�G��g�PM�_��ڥ���-����NoJ3r�j���S�冦ş�\#e��:�Z�ny�so�J_*�Z�,���t
����ߪ��T�Ya%E����T;u�s�B��׷�qq�����
�]Pu��߼�?��?��9�0,8��M�r�쩕�g��߄I�x��9 ?u+�w�S�G@E�,S� ��|JG�	�#�i��f�3-odY=��c�R�0������zӷ/��-é��щ�����G�<]�1�SC�P
U�;\lv����V�
Hb�O���<С��P=�5Q��P��@�bi�xW=���<�U������*�:��~���VZ�gb��F���Z�Ã�V�AFIO��iD_�a^y��$��Ն(/;���H�ar��ۢ�󳝡�-Q������{��Q�1@	q7�1�[O�\TN���%��n����W���I�i��j���G��Z�;�������\� Ϧ�THd��W��WD�Wr����W�p�����ԱaG��+� �vP��e�z����tK�]��Oh!w��s<t�Y�z� $��R��1`K�[�-!<N�"���׮s��r��N����@���*�Z�Ƹ���;�Jr��R�Y��".����{�] G�)�Y�&�3�ݣ��\���y�I���l�j;X�K�_`АǏZ7��S���%ɪ@|ו&Y}����T-�>�*����#��t��jԄ�2(��<h�pj�j~ew�<�X��N�Ը{��A�?���N������rzs�\��]�.ݽŮ��� ��ĎY�@ދ���=d�dV�DB�w"E�x�;��b�m�>��Ȕ�wk�����\<\V������e�8��+9ۀ�]1 �>`.5Bvc�yz��t��(����� �/�oB=׬��K�z�DH���!-��d e����H�q��KK�^nw�8(8�D jM��MU����UKݴZf���}GCY��oDmq�F�+諚�">��$E5@猞�̇:���V T&�s&1 ��2��Ͻr �;�wd�o�<��x��{�t�[ؙw���)�Cc�?jƣG�q����q����1�K"(1ea��?g��\�Q����e�3��_�e{]��''�j;�޺�r�3��^a�o�$׋��A�L'�������@��j��M�	�&f=�g��A�2��c�21��<f�,�݊G��_�R��evå���5��<`�� �b��]�u��[�E��$�Ý��48j�ӌˇ	ر��x�&a��2��?fղQ��� d.M��tE���*��#��>ޅ�Z�\�3p��cVՀ�o�� �	���X�Do����i�W�,+&̮toڹ�f���hC��8�dBT�D���UbP���t;Hέ%́l)"V;���NTH#�`qHgݼXT�P�9b�L��Ru�3�&�-X�*���R��|W y�fG6��A����vD�.��wa�#"o���P��`�G�Eq���\7^q(�2�l:�m�"H��S�[��g��u�;�񅽉�� �,���t��D�E����tMrk����q��F J�_��p�8Q���L�@��L�(�k=�X�4ÐA�aҡ�#����{��"[8aQ*�?��^�k�p�r
?��ަ�71T����O�o{�+AJL�hMUz��zh��`Hx���XT�;W�.JH	�2���>RR�Y6)2����b�8�
X6��(k]V:�˴١������J����˰�����E�FI#�nmӰ{��93�1��M�"��K��:v1��Y�j4R
U3�X���jى:�gN?�뾞s��Obe�SH�M`3���k��JR\�_`����d_o����GF�a #OV�K	�'�	������_7`�. ��E��@^z����:��c]rx�K��,����P
��?J]��a2Gw= ��kY�{B\/L9'����Ï�OaNx�Ն��Ʉ׻�Wl[�@�d���H���IS��k��ٕ��/B_Q½�J:�N�a(����+��fR�\��Q��� ����Շ.�@�����)�i�Y)`�'U6Z��OX�	�J�*Oj:�a���ɧ �<��.|	�1���>rPT��
�#4s7C2�H���7����b��%�V��ّ��}�z �����J }��L)dC��9m�br>
FF�N���[����?��L<�%��t�O?���@�{`i���� ����Z��2ɾF�w8�ֿzv�-dpWJe���!���^���q�q��c�Z�6�ڀ�%�JΎ�LA����dRO��Iry���&�ѭ���Q���r���ddAd�畡����0W��4�y��k:�Ķ�Y��r"�n*��C䅵�Ha�¦�C��7��Fo�<���N���9����,} ~v�I�[�f2���Yu^�����wö�J\t� o��4��R��o. m����P�w��_b��3�n��tH��ݡ���?���Fn��\��sN��8���C�v�%��������凿�����Ѣ��Hb�ݏ����LE�'���պenn-]x����/(dO�}C��e��X�O�Z[�4��@�#�Âm�T�y�Z[l�vcn�	���؇$c^du,V[�{��2ΐ��{$Ve�3&p�l�ǥ���3�� ?�۰ԃ�3.\��օ+�(���:O��,:��,e�������-^e��Zk��-��k�]�<K���i�S3�s6�|!����%�Ǿ��K�Q�-�~��4�0�Wzg�Ik��I���aZ��g2γw��R@�ĮA,������;Cw���q�\���?n��%�C�}�y��X!t�٥x�Q�SN�j��*o��D��]g��r�8ӭ�oH+f�+�
.<;d��{12?��0\m܌���]�(֏�V̗x@���?@0��,ծm�5�,�Qs��'e"�0>u���Kf.�P����\7�J;:dHk��7l%��"y|�ݩܿ��ي��l�,��Ud ��7��{�+��	'?�1��Lsi���",W[�FX^w�s��v�ƺ�嶺�,�n7��Qx:Q5c������0��[��P1� N�Y�o$4��n�yd���2��=�rm�� �S{!!>�L�$�Y��}�l��������]�aq��!�I�R��>����Z|�o�W�Xﴂ3���SSC��e�֗�]��9�D|��f���ʧ�Q󹴥,ΗS��x	r>�z����=���3��E5k�?�d�f՜�~�a'�o�H[l���9Dr���4=��*��x g���t�M����j?�z1�:���)���|�5��}}.?�����FZ(�K7�O1t��2�?��'`������O�����h˘�T%�Z� �e�ϖ���:���I��D9�,�-��'>R�G��Br�����#��X�Dh6RDp���RF^@���M�Y��CO����߼�j,]E��@�)*,���*��0���S�z�1`@ح����{ǆP쾩c C��t�ܝx�%T��<֭+]�0��7qz�q}>�+S	��\��ю�z��q�1?R��1|L��P�cK��W`0��H{?n5���`�"S3W^"��")~���UO����n;�m-C�W6��e��-�3=�p46�޿1��/��xz{հ]<�w��3�@^gY�nh�۔��ME���۬�eex��;s�>R��Uc2�c|�#��L�3�_D�n�
>����Wݵ�9�x�+�'����9��#]MC8�����\�<wq�I�|Lc�b@D�p��v�W��B�,¶��ǯ�6~e/��O=w͆��1�� L��k	��&�hS����Tyk���~)G/S8*�R3���a� 	�R-�^.�� �#�0G����Q�0���ٞ�y99�Hd��-��]���^��r��n����HV�	��B��Fy�Y��G�8͎,���q���e�k�J(A��^�_�L�uv�X]�
���@P���Knd�F+ڑ��(՞Y�W��68W�!�\�H�������,����������5�隓um� �<q[���C��d�,@M�} �S]���u��l]x��^jJJ�g��4�W�����{�mq�	���;�����I[c�T�_T� b	G��`�b2�i"p��O�E�k$��!7ʍ��
u3εRǸ$�|��:�`O�`i�SK�E,{~2�)�+C���٪v�m����l�n��Nf�C�����g�������}��fz�P ���|�1��+D��G�S�un&�~����5-#P��E�\�m
 `��;~<b]�����t5������]K����"�<�&Fc����
�郷;b)L�$D�uE[I���������I�Ӆ�7���e��3E�`�K�H9�ۅ+�z����n�y��:\�mOس�^��'H�ޅ��G7�_��&�6`P�/_��J+/�Su��M��M���;�݄J��py�����^�l�9`���F�}��[��/��Ӱ�5�YG!�W	3��nB�}�L�י�ȭ�$e�֣S��BZB�=��~�
�̥�C̍kn��G?f�Y���zt�����`��5��J!��\����Eu^�����0�TE���<&Q��!r�M)�����]azS���N�;��"��H����`�\77�#�r���3Fq�<���*ЎE7���_LŌ #�Ǹ&Wy�W�QȳԘӀ�)}[�W<�ӟ��Pm�~=JWn�$�27��+��ȳ�$7�U����N�$A]r�CSBF�&w ���T�O[Q���E��=��=�#a��NRN����B��I��8O�P���l������
c�1x�t�~jR��/�oB�c��s�҈�4�����۰p����S��l�P�h��]��s� ������6�>��O��k��y� ᫘����_q8���')?J2�|i������}%̺?n1q����f�}��K�������7�Pڗ8R��m��+_�D�b��}IFp���}��Xe�/Q�?⎙��-��X��1W��E 5��_o�vi 	~Bk���7�#�X{�RV�S����7|.z3Z^��%���~k��\���G�`�&ːPc��LA_E躂G}��b�d��Pγ���Z��g+Za�D��$LҤ�3F#�}����fܒT�����K�cc+�������q	&�����2gyC��B	&�I�g��|z#7-��;�+���l�Jy'�P��x���1-z��������I=�[]��c���3V�Z���452��k��{'C`��S_��E;���t"�(��2�t���t��HJH3t�Hw�Hww	C�t�{��{��2g��g�Zk�{fƜ`j���k�9�)�稴�fC <��{��I)h��f�g��Y�=�!g�,F�t _�6��pko��$X���b,=z"����ԯnf��R�<_�yM�<�a���z��bT�~��2Z^�h�twS�E`R	���T�����r��${6bŇ��Z�i�S[jR@(s�8G�+??�2!�7W��֋��/$��ކ��ߖ�GoP��� ֊�+wc]�i�.��5���q&�b�e_��d��"'�i7��:B �-��H�@�P�_0t�0 �J�����	�s�lwu�6<>����v~��8M�{��'J]Y�.��_�Kw#�C�?�oai9�U9����"4^");��ݝ�~�b'UN��	�ĕ��<��)�m��0X����$H{u�\��������
d��Bw�QF�6��V��>�Rw����Y�\a����=��l�ͤE!��Wn��ڵ�`�1#��k�1�y��cP����&�����Fy��n_�����4HKF ��VC=�K�np>L���j9�ȩ"5�C/�6Ө����0��Ð��p&�f�S*!�ک���Њ��ϖzE������E Mv\��MĴk����+t����$����]��7ֆ�S�U�9��c�6��xG��|'\Ѝ*=(�u{'C`�Uk��~Q;���=�t?���D�x�ǻ�T<�{ƭ{S�5�1��ce����D��|n�k�rQ��Qn����/	�`E!`ŔV#Λ R�@����v�����O5���P�p���Ȅ@\���V�7���o�YJV���I����l��8Ј�\f.�Q%�6|����u	{�Gn�n�r����g~
u����呥���f���M��1)ۂ���o�V#��W�0����ߢ�}��^�L+t��54��/��xA",ŗ������f��o�+�<��^}�W������2 ��|}�e��L���l�Kh#&�7����6�����O\G�#d�'`�ԋ��ZG�G�&+X�����8��;�M�.`E��A.q[�&�Oj��E�[Nw��^%,��j(A��-&�,��,P�j���83T��4��C9y<u�'�C�'.�$�XM�����g�2�|�N��Ab�Ƶ:7Tmł�$��dy�u�˒�L���<?�o�K��ƭw~�	�O`G|Ά��g+k�k��ۚ��E��/��쬔��s��CYڣ�E�_����a����nS��Ae��2���	b�6�n0��-k�r��HT�bɤ����aθ�j�%BI�Zp����C�:��(��~��T���뼏Y��@��
��,��pqk���� 3	�r�������D9�{fʴ�#�Z�K'yU�h7�_�hR���k�H��_s��ǜ,�+��k>�B��~��A/��ԩ)�$>t�,YxK���}�z?��E�ӃIinp%�J�c��{�t�G.��kcy��3e�A�|�!��� J,�կ+ތ�Q=�`W��@:�z����y���\�]�9�~N���m�ڪ�N�*OEA3�Y��;��o#���H�S�|׀ד\������-T�4;�Ş�`~��e��FZXN&���Z���%'�S���+l�g���=����t�<��G]�B�dA
��/��>�h��4Acz��Nr~��=�g||u�^��g��?`��P���������#��i��x����qCU��U0r�\��U���tq��xəf���^btH@�u{�t"�%��5��?9����<��fW�l��R�����7dT���+!ұ?�%���>� ��j��0]�ei���أ%��r&�|�Fք��H�mO�� ٹ��w���?�]�&����$Oa@	J��O��r\2V�X:&��(�����i�5��K犯7ʍ�Q��D�
k�k�z�k�_Y��kW�%����r�aap���'jȈ�Y�噁���<oW�H��7�nk���b�=t�S�h��Q]�����VE�t�V�Y�s	y�P.�t��q����@�Oy�'�b�V��o87=�'3\�
�5�'���[�u��M|O�uV���|r�Өx�}y�C����g��ڐt��!��cŞi[����9�ᴯ�k�`�rS��I<',/�d6��6WP:3����Jz1W	��`p�L�v^XX��SN�V�)�!�&�f[��ezC�T���3'�`6%)����^�eQ��	']q���X�Ǥ��O�Yu`qsT�����\�12&�=?^�i`�QW��=��3�C^��Wi/��QbKmϞ�S�n~�g�s��=>���?t.A�CiX8�t��Y�h�|���n�����ᓸk�{����H��O}Լ�{j�GU;O����-�30���g�gW����^�N�"3#hW�|�~�
�H�Z��s����(]��{��ǖKY[+�Su�p3F��<��A@�����=��3�����D�t5N��b��6�Nc�~�d�N���h��g��u�����}r��xNJ���v=j{0���7�u|���D���P��q�.|}�j�L9�������
�_�jb�'F�$W������oŞƩ�q��mw�� ��.���8�����]�Ac�eT����	��Z��GSl�s�r��%������lug[�Z�N�����%l���I����gb���h%�n���D�=��y.~��W��<��#=��#!��q��&��n{�l �_S���1O����]򬞚���O/5���[��o�*�V!Y�E�x���%�=��o-;�6�VD �=��n��œ�fH�&����z�$_��Fosf��ص��I\j�4*�C��������\���E��&)� ��bvCds�zj)��WD�k	^I~���ye7�
�:ś�[ݎk�H��%��Q�^8c��� 3������5V�'b��9`,���#��3��[ޤ�5���҃ˏ�/N�g���U��kE��b�F��)�e�D�$y+,8QVo/�~�a��ۀ����E��Gz(��{�B��"('A�����^����d#���R�g�j��D�"�i/����V�9�4����D5,�o�< �|��F�� �!��H/�aO#�&$QiMe���*;�&C����a�oJ�	]��K����q�^��2�B7E������J���Q(����y76��3����y2�f�\ ���#�V�Y�]9zN��g#�k��06&g�z~Q�o���P1ٸ߆��Q��}	�:�wQ���1&���(���$������}I����K�X��KFQ���W[b�O�볯��?���F��<&a�喞�]"U�a�I�&�L��`	�$�=�Y|jڪ�|D�������{�zǳJGT3�'� Ւi;V�ƚ�X�� )��9���<�z���2���9��a9���#�C�5m8�35R?d���1���j8�ga�!QP��Ѵ�!&tk:�*���8�al���n��I��~�9<����mq����վ�ϵ\�z�C�8�HH�s�`�E!m�mB�����1�����@cT+	�O���30 ô�q��P�Ȫ��ﲥ�&}CN����|2D��l�?M�]n���h��k�2@Ȣ�W������rm{O ٚ�0�'/���R0��*8�3��WE�m�zJ������7EX�?7��g{���ҙ}��4����%Xu]Sy��ԡ��P��`0�9�_~��}&֟#OS��>��񸯤�{��ዶy^ZE�D�1z���e�>v�E�P9�
y��xg�ys|1+nw;����^$����7�}7��2��0�������Ͽ
W��Hٺfi�E�9���Y��2.�}5Y�T��־�P�y�����>�;������o��;o�G���i@"��3�Pl�1�9>���Ԉ�ܮ��3�b�,�>?����ҟͨ[h	�v��0ۏ��HR����He���檌l*O7:��]�R�u?�9�} ��r8�tչ�d�~��x]��Wө�x%�-_m)�|�C�����9�$m�Q^Pa�*���%�����I������qɣ͊Co�³����]����p[����D����|��$$�ҭV�|������w%���:c�25/��@<ёF=�:��j�c:#�Q0�����a��H��_-����!�ji�-�j'����?�����d�wݥ�������l;�j��[��oa�˼����:�Il���d_%in9y8J����Js����9ʠG��pX*�s���y�!���IL
��}�4�r#_@kh�L�����V��$_B��+���62���t��n���������2��l!���bx�I�z�H��n�_���M���/�)��*��Bٓ��渼�ʯi��J{{�[�[��r���M��n��?bO��A����VA.�"��wy��g�d������{�HYf����a��U˧�ǒ.VJ���~G�4�w����G�ڏU?��{bv0k}%ګ��#
	����(/�r�]�_)�?�,��>���ϣEdf<�қ���0es!����U�.�M�Q�)��]^9k�b��L�6X�zU4�r�� ���?[��X�|k��2w��ɟ���~�IC.�#��7v���Jq�WvT悥�
�घC��
�'kT�-Ё����E���,�ݓx�gg�t������Y���i��oB��efi  �����蹬t���R�-+��NՏ#�
s����=����ܸ�;P6d��YNVrhĈPI���pO���Kvc�Ȥ�UX&�w@_s����p�{^ׁ�H�H2N����C��ēƔb�z.��f��F�N��z�\n�'�CJ���3��s��ݭ�����Lv�Ή�h��q��y	���=l��K+AKn��2!p���jn�� �@Dx]�d}_Y-u��m��2��Z��Qǵ멟��eM v˩�����*��͉���(v�y �6��Zf� �r+��:wk�+��
B������t��%�U����Ђȹe�W�C x�'k3�kXJ
D�ii 7�%@eg���ʥ�
�!n�;�0\��!�$OF������{��N�7/�ޫ���A�H�3`٩�BG��M�����
&9���l��ZG�	hlm1z|����/Un�Ԯ�Y��ݝ߸�p�8Q/P"jg2픛�5���f63��:��7-�n����B.�k�9�\�u�d77�8coz�[뚨hWC�VU1Ӎ�bdv���U����WTHFw]#�`�/�����N�ߤe3���>[;L��ai�R�?�����������ۣ^&�琗��笫�DT��=Y��2jz�&N���H3i�=�'M�.q�����$�$Q����:;w�&ߴT��j�kM��Kz�Ǹ5"a�ܬ@94"pg׳������OK���wA��5�B�x�rX7J ���!g����&A���I�i���|�{M�a��\��H�Z�<gd8����ϻ4 �w�J���-�߾[�P%�@H�ۈQ䘶�GD��v������D�����e2��3������Y%H�)%��a0�yTwr&S�76 \z<���
U����xt4���O��C7Bؠ6w�Z��?���[ֱkw�{�G�����o+׆��뀠�������!���/�C`}:, �v*��Έ���D���h>�c]Nt��(H��,�ͰO���Ԙ�ID�n.4��՟��[��C<[}P�^���ӈ�� �:��+m>!q��$�v�U��C��#���si�?�����o<�ˢ���)��\�/t�ux�f}��ֹ{�I�@�Q!'Hj�F�
[��M�>�q��/Ƚ!-Y��[���]�o�z���,���aj��QȻ��m���|;c_���@R����/ϟ甐��4 ��F0��À��,��p�/{S�L��8X$�?u�~����5CQNN˨ڴ�p5�bx�3�='����K�Xx$�0N�G[9��¬S"��~�\+�<�R�c�x��; �>�(`��66��9ڱ(���'S>�q4Oc��eN�,�f�w.�gy������z�6���~#9��Bɬ12�Mͦ���*]%�E��h�;E{A����cBnɻ6�fGϰ*Q	i �F[�?=�8F�-�	;���]�_��h������n���I�O���Pp���ogT+�~�����ݺ�e
�L�^M!�.�"���)��5��q-�qG��$��hL���<�A�H���3�a֨�R�>\����3����nz��,��E��,#�^t�=u�, �!T��m#F���@f�]�;��*pd�F2s�{�x��"�2Zf�g����Q�|�v���IuN{y�Ϙ'�Ȟ��?M ۑO�5C������2^�aJ*��vߠ�Jh*[�P��Y���������A�#�k�t�ce��2�R�� ވ�;���� HUx8Gwq�]���W׋�vL��9��NU�T�f/l�u��u����Ң�jG�]���KG�-e��r�?F��;�5���W���B��5X����[��b�x��?r�l��kG��䦖���çi��74�0�U��C�\�?�F�h�k&b^���S
 � ]�Ǹo���~r��@������ D��׮��5��t=�洘��Y{c�U�b	�apnmE>�F�c"�}M�Z2�WU]鑫�*$ �A ~w�X���ujr������j� w
�|�֠~{�m�H٠�<o�h>�g���Ex��j|(ݖp�]��4�������ϸ�Y�1n�}�T�)]k��Z(-!�@LmR��~f�/oHٗ;�B�&NϹ��U(^���xY���kV��Eer��X���� f�m��xAz��e�AW��W`��Ů�́ـ����c/�2�Й�>1��K�z2�6� �D�uj�sg�n1�o�%6��8��ZWo��̏�*��'
�>��͊�RՀPwT/ZOF��8�,�|��@��Xh��6�K���CR�#���h�[sdFĻg� ��(���^4�� p�z��z���8�R۵7?�!ꯡV���@@�n>/�!!�O������И�C�K���[K��<�3�"�TOc>�����iql	m�oo=�j����|��pė{@W T?�����A��� /<a�	Xp�G�d���X�E-�"b��G�䂊
��:�����~w%�q7����6���"v�~�,Jr�j}�#���;L�V��q��2��q���Q߽Kb����i{�Q��@4u�z�����'��'*���ATYy�vp�M �*��e�,��H0QZ�Xu�!Bg?�@R���2�X6\�(/��k����B,�j1R�N�$7o?j:���Wxq�&F`�7�y՜��]��Fy!�2�ڃ���@��y�oot�_��?( �������yt�F����3�6�4��f�O�����A�h��,���:Vj@�A���Y�f��Ϭ���y����l�h4���uX��s�����n1[-�jA�l�"�r �rwG�I@��I$r^����&ށ���~���EJ��Aa-9�ÄV*]7�q:�}��N��v4(G!P9�B6n;������x�mzȪiIp7��Z~�OT)ڜ�3�uʔ�6<s�w<g�:���x�"n��0����7��u����-5Ek�d��]���ˣӌn��h��Ϥ-,(iSt����%��������ap�˻��el�2o�����@��it�/��w3<��F9!
���%��n��@a@�:@���R����R�<�yڀ�k�\:3��@k�<̰��A�����rǤ�374��~q��z��8e�"�F�vG��݇0P�~��
�$��THI�S��"8���4F�� ��rk6�I�v�S�ӨC�j`��/P������nO����$rs�p�>?(��%�:�w��6�8P����/��L}�;�#I�L�w��L؞���<�D��i����|�T�,�ż�M�nh�g\"y�4�b�G�%F!"��g���\��	�/,����6Sx��\c����`3,Z�َ҅�iTl�#7BT3�q�DUm��Y+
	�bF��U�0�0�5((t���w�`x�p/KG`�����S�W�-��/��YG'���L�������^y@���fk�".Nw���{З�j}ܺ41�Y}4����㍫������x��V�����8�~[T���d��o�f�cB��ܲ�}���-c	�b�ka%?4�������󭍏�і��@�l>R��&��t)ǯOh�!�&���2�0�� �N�������`:��?���p;��0�0;�����Z���u�?�_�BL0���f�v�_���OM��\%$ȳ�S�zQj�<�sA�ę���ֵ3���|�r�1,��@%���'\��6ʟT����?m���3��ښ,ѷb�q��^�AǎARmv�_L�O�ne���nn�B䚍����C��q�= ��#ϔ�6��������C1c�F�R�	R1����e%G�V�H�)���GSd�h�5�3H�n�|z�5�kC���E��C�='����h�v�w�K�r�o��)0c���"�ΰ�T�|���`(����\2�%�vڍˮ/���W@�L�?�|�h>9����:��ׇ�]�G%����.��x�6_�H�����Y��&b�Ƴ�@��)*i�T���j
鑈�O���<}Y�>[X uL�<�Hr�o�|�i��|LƢyO+��ɜ�]:f���^����kGwzY��_�I|( �۶�w��j@���їvRc<�l�ltk�)_���t'7��.9�;������^ߛ}����+;�zP5�LJ ����>|b��R�h��,��v��4r#t�a%Q���� �X�qGڼ~��Yj���DR��i+�41�MQ�t��٨#ԕ��>jO�Yw�#I.Pg�u%*����{����L�ȈQ!�و�����;j�ӌ9���8Dߚ�,��j�BҖ�ܺv+X �B�1_Z}�[vvs"&:J�h�����r/RQK���UNA�3 ;Z���o��lL쉏eJ2^�zO=�,�5�{j���%����� N�����O�4��{�&�؋��q�@l�#/���DNw����>��%�T�=�u��g�6N�4��f B1��"Gv���*	�瀣A�Ayj�� M&g!�;{Φ��i�F9���������|������X�f�z%�2�(<( pʌL�pt����w�*��H?{��V�=�5V@z!t�Kz�]�a$���1�[x�v�q�w��EA��AH$�=��B����N�s�)��(-^��;���^�_ qG;��a�𭨤i���[?�^`�D�a~mW�o���9�c#W����P��7�f���E5�ʍm��{��P>�xg/�ӂ?+?���%��T�|q4v�������]�x��.crܙz��5Y����sUG+:M�k7�����5�x��ʯ��:���	���ܕ���ԣ���� u,-S������V���6�C%��&��@"�-�X�[��'z���O�`�$7�:{1��zNRAΪٷ�&��Iy��]AoX��d0=�ϩ&2�p�EVU��u��Kнy7f9�vU�g{��ƑJ�,�����:��N~*d�<N�RW���{���~A�o�ΐ��y9��Y�UCE�ج���a{	�c`��x�F��?F\#�@Jޗ���X�)o��v���L����'�q���u���>�n�N���)^��q�TAYh.��l2�Iz)
Q�${n_Tv�Q��+�ϊ)��y~���Q��$v�.�uȾ����%Ewy��/�a)> ��լ�l��z(��oTb℁��1� ����qT-�����Hv�%W %d�zg�2����bV��x�Ǜ�O��ú�NR��h�<�[p%Um�
#��h'P��'������l?�GP(x�i�A�T[F�	�*����u_C�D:E���ߏ�Ph�y+0�q����ְl�o�!������V���s���M6ӛ���[��ꋣ=��^#��3�$�F�s_�����x�5<��z$�I�P���8CG��n��s��9���TLX�.�硁�'L6��eN~#���u�	�91��-�.���\0Ӷ_ǥ���x�9�ůhH��<�A����m�H��p�8:B��p�hۣ�=��^o
�⿸���[���.x�-�Qq7�K���r����3��Ѩ�S��zz��.3>t�/eZ�u�م��خLI@���p!�F��6�Z���K4Odx O=���t���=�<`�|O����1�ln�	��U� d/���a�D.�A���^)�D���ɰ�����9��Gdi�#���}g�ʼ��9΁ȹ� ��	K79�u�R0}�D�2h���X�H,�Z��a ���A�3PzR�&��v�y�G�y��mEM�z�q�zLpX=�~���ћT��}B� ��+�<]u��}5������8�i���{�g��Y�k{�����)2~�摶5�� �H$�:�)!�ҝ�S�ed���=
��x�J����"O3K�D3;v�M�� ;�ϳ�^0\:48��LvV�c���$������[۫�GW���[ �/����B�]��~E�SZ��t1	�稟�m�﬜����̛q47����oZ����5���y�f1}2p�������j��a�T�(��)?�E�oԢۤ�3<R[zK'lID6�CI��
F�$���%,Ny�~xT�[��&�6MRV��N�H��i\~W�3��~�'��� I��8񇔔Ժ�_MH���9�]��� :%%'��2_�Z���)�a|Lֺx6�h�->�,X3^�߲*
=S���ix]����a�ZI�CP�i^n����?�����3>��c�H����N�c})X7�+d��6�	���Z{�9��%�����\�(��JG42Q|w�aJ=����`ũ�B�ˣ���Fv����+��	�W3���G��ОQk�W��R޾7��h4ߕ�xf�m\C!�m���-��|�YuP%�V�0|/Z�����O��U��^8��d�����3jb���ڇe�p9�c���n	����D+�C�lF�|����&W����f�J�=o���4���z	D�)�VZ]t�C���-��;uƮ���;q �^}�2m9J܊���>Y��9� �A[�a*�H6@š2��V)�(4�zr2u_�1�����x>j��y��}�t��ʣ����u�9�1���A��o�X�|9~��1�'���fQ�P�Q�z<z�O�P���YWz=�/;A��z�/�<�hi��I�1W�y�:�w�Ŀ�o����ٽ��LoԚuj�t�_Wy��ئg[��X�6�<C�D� ����l��*I�� 'a��ʝS�v��/���P *ވ*����.��o����;�D�1D��_���늗�+Ƴ�^����n�2Mڀ�}|�3�]��")�Z�����7�u����ޕ�=0[��W%1�&n�!������c�cV8Z�����:s����Y��!ro��or)X��(`N�o��0�Y&Of��MZ�qN�C�������m,G�w4�Q���	���!Gs>�3ݓ=~��76�g�s��И�=�U��o���Ã��5ї�L��E���tܧy� &��=��`����F��5^v�����n�(^��1TK�F��o�}��#u����*����ArϩQ!oȩG�.�I�j ؘ�8��u)��Wɂ��D0<��Tڋ<�Z�0w��8��].W,��}�X��um��Ǵ�֑i��Fe^^\
U��?&�
H����4b������-?�")�N��b����R���o�����{�1������z
FW���x�䠉m�J�#߫bI4�ɢ���f�
	�ZgS�5�|Q�~5�%��=M�Eju�W�b.,��]%��:�w��i�!�8��y�f�D�-@��y�l2L�J�~�M�p������Qȕ����� .��8���@�3@zA�-"Хğn�XH�m\u4�Q����*�a]�Ml�ʇ�Z�\<��������6K�Ʀ�+%�P�S`��&?;J���S��d�u����m�J����qO���b��b4B
۟ �� ��ܛ��z������3�����h��0��[#��K�E2���B;�����|wޗRr{|�~�ۑ9�z��3Ƭ����#���~|�v]�o�hb&�IE�{?��D"��aE����`mf߂y+��ލu��S�ʵ�}5kņ}=�Phd�N#��Ff���Ov�ٜ�ͧ��G�Y�?R��f��N;,���(<pܚ���kr�z�Z����?����Y��M ��f�Q���&��� �U9���'� /�qj#�h((K&I�V G��n�vm���S��}���hWME��9ޠa  |a'p��>kR�.��O���t�.�>>���D1��m'���Z�]��?��B�͵�܁���at$M�7'�����2��*��9.xsnF��Pa�'+��7�"T8=��裨/ˎO2��u`��fs#���8SSa���6����.w���	}����f���eg���$\L4��a΅��m����*�z�>���=�n���*J"+���)d��M����U`P�zb�>��v��~����ʺ�}��>}�A�⛑c���{�E����w�M"���/�X�v�_�Y�U���s���Wˋ�
�u:(��&���q�K7�n˒�^���fdVEţg<�! dd@ί=e>;�b``�U��yٱz���'�ms���%7>>$P�-�f���j�gF�>��\�/�C椊���t�YC5 ��7e�6��m<��W�&eߝ���<�'���m�����i�4(�C}"jj>���/>h�Z�:�n='[M��ų�Jp�n�,�*���f�scʋJ��<m�x�re��]�x�X��!���!�5c�=��@x�����_��`��Rsm��S���޵;s��%[�f��� J���aK6�@A���=�,�����6p�%��yX�s:���}0cN����O�7--
�ccszT�@u�q�P�����ٴ�,gF�߳���S��Q�6�G�[p(J5���ȳ�9m˾�d�\��y��ܗ�.[��)M#+��Gр),<]c�����e����U�(t�mJ����}�ŧ���<ER[����p��Os�1�c/����Xm��=CW��Ã�P�5�^l<ؙu~�.|��<#:/����P����8����fQtgk��gv����D���8�������`�Hj1�lqnZN�ZR�1W�Zm���"��|I"!�N]P�E�OY4��~��b�2�!�?E���ֺ�H�2 3X��ރ�����贸
2�����l���d(�8��2��O�q�G�_���m�:B�/GT=�fYH�n��o1����(v�O���Ne2��	v�Ǟ�er�@n��Y�;JH	BI}2�ҢikPwk ��?���S�P�	s��!|�u���wn�;<�KI�
��?��i0��-%X�vM:��������?��<���z<��D��퍎��9:�ܴ�l�;�SfI�D���F���L�v��a|8�K,�:��iWZ�K�o�`V�Kf��h��%�qJ����"����~��:Ӕ�.+kC��\��A�i[*��*\8��BE�0�}&� Z;��֝�UTa������� �_hɔ�08��P��1&.ePT���Y���O�wr�)�OҥY�KR�RRe`^�( �2g)�;�f/��$��O��^L�W!h&H��� 煐(�Z���}4���rS��K��`�	���x�"�DCq/v�~�02_U�G,�Ѫ�YN`���ak!BJ#���)�Rt;������k]�������Y^:>�fX �h���t|��s5ش<沈8e�8��rP����K�O=Iϖ�85.�3�.t�i�	�<��������v���CƖ��/�~�e��gu��̜�#��Y�<��d��Zz킺]����)�3̇$[��3k;_����Y���!J�Q�K5O1��M��q�e3v��U�>��8���-��yGn�uN�D��υ�E`8�
��dj�8�F/x�:nAoJʟ�Ҏ䘒�.�:��Ƈ�c5�jh����X��q��'ץ. c�K�?� ��b�����95%#n��j-	u��V�Ұ�+Q�g��T���|kiA��>�5�ʆ��O�|��s~c몕H����<��4|I��8ʓZ���=s��t�G�	�L	�z�%�$��ᠷ��K6t���;���M"^����s�Θ����]�ͥ�?�����qfY_�u��=�b.!~$O����Bo��!7��hW� �p�l��
l.#1z�"�G���)"�6�s
��"U![���{=5���eUyR�r�?��+U��h��DB�!<���a�|���/x���v%����X�[u�U���N����U#�z�e��'�+!Ƹ���9��XA���ގ�*���}���W��D�5�:q杒#�q�Φ&ӃY����/I��@��[��c+�05�tOM���q�y���i8��	+|@�߮	��	f���)"��kkk�-�/�M�ab�@MpX~x��t�$z�(�G�f�g�棌�(}�Îu9���$L��>f����9E������S�cO<��t��"�(�S��s}ˉȥ#ɺ�`�����U%J�y�#o�Mʃ� �R@���:�R&5�<�z����麬hO]u��$�oK"�����3��c��k�%������1yb�*�G�CWBA���w��z���=o)suu���ZHu'��٫olw��Kٶ�-��o2��E)�����~�v0���;S��ym%4Qc�Œ?r�m��|��ӭ�|!$!�����7�n
�?"�z���,�!���!.$��$���j�.�J�uix8��@�_GLœޡwI�,v�,Z\/vD`��O4"N׃$�Iv��sLw��0��C��?�4�� ������̺be�r����y s����)$M���1%��y6��BPa�;a�}������a�ү�J�^�`��E�#p����z���V�76�̱9T5�\���6��0{��e��H��5E�ddM3�b��F���ri���>��B,�ⰍF��	�������[�^�:c����E9�:�kq�h��r?ry���� �Ϊ�/tl:�5��&�)�`��F�o��9�bq��p������ jT@���ø_q��͘�9�&�\������]�3��Ƞ�����HI��xC,x�x��!P���#�y{'!�~^���Q����<Z��*��;�r�_���t�Qci}V�����˞P�(쀘_s����=K�~��Z)����Q7���RI�����;�+!�9=�	p>߆�BZ�.��ׅ�eo+��n��d���F�U��:�.�11��w�;����~x4?�AT�u.�5��ف>i�aI����ヂ�h��sa[%�t�r�H[��W�]�%	�m����Vb��$�&a(�UTw���e�Urn8��
<}Ϛ�6)!5������%�&o7�%��;�;s|Q]%�C^Ĭ�U�f��;F����zؾ���#�v3�42n� 9�q)đ6��(�0��Wp�;��&l�|������*�<�y^�1 �,�蠗4�������7)��p�9�w��B)5���c��0j_@��(��V��ńu��� 8/�)
����YT���y$)��KM=�mMz��r�B�V�\tDI����<%��i'��@�V�y檜���z��a2�"�.~�<��aS�,n�Z<=����PE��vƶ��dd��o�"�L�蛏i���]=J��>2f��	6���W�;�_<�ij���۬�XsrB�F�m���Q׃����-�������xϋ�c!# �[��O�k��!�^�W�[A���.�":ۃF�� �+�*�~Kr����
���.J��ˀ>\�4�����,�I.D0^ `Tߌ~�DR��%��)pǭ��T}&{�ܶ����؄�&���ڐ"�k�_&8�x%��#�:s�Q$�h�i�k���CV�QC�K����S��m:U훖�jd��<ajƭ����!fneݜF�定�15�'�'�bǔ���)� >����P/������#m��_�;���L�j�I.2ԭ`̟lO��3{<@EMM���r�xF{N���:��՚q���-!�����9��M�~+%�T�W=||�쪝< ��m�_7�̲�e!���а��}S��F��A�B	� ���R�����)��du3��2�yw�֞9ק$��weh�]>Q��[��Lx���{�Fg��An�Up�I�O���h����a�����'ĤHv�}�t��U�f+�sƐz������2�-�vs9�)� �
��O
������*0|ȒH:e9��E!q.c�?��P�\��0�����"7�U`p �f�p�9��t�?L�갟��.C+�u��,���b�cKG��.6�U���9�W�/�6X*���k�4�NL�B%z]=�p�a�Id�[�f��;��J��"�.�$�'��f�:pUsW?�ޑ�N� �|Mn&�ZuO��z,ӵU�	q����:j�aB�G���&�=��^�n�$AM�ğ���i��Ȁ���gql7^�%)�n`�o��H�=�(�wCė���=_yW7�����H9�C���Er#$"����Ԋ����i(�X��6��o�l���Ё=��zf�1���r,L����*���Č�r��L<(U��/S[��>�>q�QI��V%va�}�SKF꛾��$��G���CZ#�(�=\zNX�w�dε7[B5�1�=`��@:�

=�)${/����
���7SU[ܽ�%��W:�g���A��?.�P�����}��o��#]����+�7���)�t�c�*�c��t�)��4[ZE#�2�ƚ�]���4P�Wc6���](;��^���~~ÿY���0-���{�aA�Cqȃ�Sψ��z���.lXDA@@���S�[�D�D�d`hP@J@@��n�����c��?��|����֚5�a�����}]׾��>\�u��Z���Vu�T��u�8������!���+/�������j'ea<���NKuN���S�#7=�̲��V� ��		�C-p<�ʒފ�B��?�aG3hb��������U�=_��}����P�l*!,W��#
$�,o���i@B����L=I�٘�V5_�ϫYU�Ze��*s{�rCq��3���R�gdCKcfw���//VA~�˿i�9�!��>��qc~ dJ�y?��]���U�&������I$�-�@x��[6S��Z6�:cTTԄ���BlJ�(��ar(Z~�*q�rvF�j�a=�4�;X�xxYJ��k��2�V.�,J�$���fDE�$N�.�$��DP;�hŵ3�/~}<�:�ɱ���LgX�}�;&��$��l�+"�\��Q8�.���K�k:[��#>����$�O��R��Mk�������D�A�뫍��!F�H��*��8x�cԂW�x .���y_��GלU����恟f�C'*�g��˽�����=l��C��B����ؼ��l��`�L�& r?�	�S�s$�\k�$�m5S��pui�Io7�˙�5TW��v�&�J�������LE�斥Mf��?^�n���p�]�9��<�V�<8?	+ϧ�ST�U����J��Q��vf�*�Wܒ�P�zȅ��������� :!��i|�p��hy��Z�5��=a1�<_������>k��,�⿄��|o�������N&�z��N��ʯ)�D��L���tq�ϐ^7�^Z���;�u�ퟑFsv�ݯ񪟪\��"����/����hꡖ���'�g���
)|����z������UB ��\<�-�����oa�0�q���U
�m����X�}�d39qo7;�acIr�����X���{����1��]�D�'B�qٗåa�73�C�b`�`���D����~mǡ��������̠vT�YK��t��5S�&Q�K��q��}Z���s'�I��t#=.(���N'�A+�X��S�٩�Sφ%a���F4.>K\�g���˧Uj,'z�1B�H�Ȇ���ug�I|L��G�R��k�{G?�  ꝶD�����ձ�9�ޓ- �]) #��\T:��	�oϮmG��O���.4����8�1����NS�d�:���[��Y�E7�v
�c�ц��,����B��;�/�[W�8�G�;�:Ri��l\%�KRa����w��4x	p4�&q�֭�U����
$)*����6�Ӎ;5�� ��do�94؇9y���q�^��e}�^C�q�f�����E$\T�^
��y�I���̢�gf.*�韇\�vX�a�/!`��J���
�:1� �2+ţ��2�C��znNO�y��s�kf8������H	Z��裫�	��Q̣�=���UU�&~9��	`/�u�h���ck�]���N���-�xA�Q�d�ϒ�	���z{T���Lu�V�pE�ֿrV���ok�!e���Ob#��_�����v�!A�M_w.��	�8�3枙%g��C����m�-�cF�dN(�\?M��7D=�@�e;'��
V���a����`�7�Z��%O��i��{�qv�L�H�1� ǌ>����-�'|�XۣϿZ&L�k��@�ud�ݚ�0 ?�08��W��3�Hw"��6tUM�@V�By�/)D9B��ab��<�*�[�.0� �� �'aM���&�z��K��L�L�VxVh�N*��vŔ?�����m�󥹐o؊��{�'�'������]�O�������w��%}�v����j�l ՝��)� �n�uE��r�ߑ��?nK�Ӣ����Z�a��_�46�@�dr�hS&��:/�D)܆i������O3����CwIy�89�MSe'h�+����*v�������I��@�')j�^���gڴq�`����bҡ�ݩ���K����a|D�(֋d1�7	���a�* �j��DM���l��Av�D	OI~��r��>/���JbA�5�W�ܔ�gA�@J����4�S2�7��YQ�ӝ��LaJ�*g�g��~4?Z$.�U��|�`��{͇%'���U/��>�W�v�?���T�`�ZH�H"Lh�T=����Y��e��f,��VWL��(���9:ύ{��5�n����j�3������M�W��(�	�ff�te*�z�e������Wh�C7�CPz�{�D�+���׾1A��`n�"��[��<Jsח���xw�/�X�r�IU��4�i���N�8#'\W�J^9Y��1FK�Z��<�7�P\e.>,��g�a��?��M��I%���cv�|^����,����%���T��#a'����ka�{��~���s���Rf�K�����J?��q��#��
¥e������!��x��eg����8��LW�.W�(	�FU��5��3�K���*`Y�g���޵�J	湸��>��ez@X=1��>n�����Zŀ�0�ڃh���?�e����, �^���u�Չ/F�(���i�q �MO*Ĵ���2�r�j���j�@���
�}��k��� &�ﲷyr�KI{T�M�Rg>+��y�C�)'�Ѽ;Odǉ��LN���m�P"�D��a���X�ϲ#�tZ�	E�c6�%��w��?Y�R?�k�����G�����`uv�e+���8T�-7eV���,�K�R���c��$#��)Y�L:��m��NK�#�f���k�;G,Օ��*�o'���29HԶ��^�@>��\�)����N���#yW240R�'k�B����ym��ƟqJ�+��?����-�_�,6��]��>�����3�Z;:[b�~������aWr�t3�=��r&����ԋo�Rj���ݥ}���4��¾/ofo�D��G�|n�l
�a[Ź��ݬv�7��x.f7�vȢO����LU��K�	STL�dmfA�C��+rȖO<�*����l-:���c�f�%�QPb�0�}���fZ��F%����}3h��V��K0�t;%�-L;�E��� JM�M�4࿧4@��h8���Iq�?��ɑd�������!��;���3��o��r�Ӱ�!�cMr�.b^R0�;m��q`���~Ba�,[�g��JKѸ'�̺8�
�7�����m��p�w)��?E�ΌÍn�p�>-�����|��[֧�@�W�xJY��q���z����F�WX�@�Ym�e582�J��s�7��{�y���*q� ~vQv#�li����b�7�K
,�abwW^(�D>L�������������u� ճ���Ez;�F[�K�1F+�4b2��iiAU,ݹϧs�.���F)�1�
�x[a Uя_H0��+p�@�/������N�[/x�����
Z�ֻH�@�8�o� /Ltw�C���ծH�M)�����'�:�	�$��d�/�3 �H7� 4D�vTQs�M9��Hs���2�z_i�-�gFb!���d��O��2��P����=}�z�oFh�b�]2�ﾪf.	93�>�����b(y�ғ�*,�RF}sв�>������-�{Rϻ�-�#ذf(�}d�2&ל�s3��_�D�����K�%���y�A2<z,�o�1�D����Y�/e�eA2<db�=�gu����|�οظq������T��/.�E4�֔1v�kiV��eD�I_�� ���A�M��p���"�'��-��*����Y�d���N�� K�3���ܾI�i��v鰏%>�Z_���?19<���!,��㲜@���y�s���
M#F��7��_��2�+�NT�͉��8*�5s�ι�}+f�0�r�R>���-��������D]*O1�F��f�Fj	�I{_��A�C5���\��ɭ˴߮�w~�֕J>Oؤ�>1��%��<e�4��O���?+��tV��c����� Տ[}������YC�e���}�T�W�n,��w�AmR�j���<����Iҗ�A��=D�G:�a�a�c����Nʧ�=���l�a$�!�����Y�L%�8� �O}�Â>�+:�F3L^収?;��ev��H���_=��Ind�O�mr^�v=s1�뫰��p-��M�Xő%�F�t��y׃cY��aY��O�}��� �E6b�G����A�5�d� A����M�_�fw�2R�9�_Kk�{�:���5Y�������U��R��!y%^
@��36���6y42��̃v�(JU�l�[0���B�5���y�R�G������)տ�,�?�GXZ��4�G��|�촌��������!3#���p����A����],y܏ |���Z�G)Dg+��͔r�1��gvw��ر�G�unu�D�B��������hƊU���`J�J2<�؛U�9���]*�Q]�sw1Ox�|�����tSm��Ʊ�,���
�3��a�Ȗ�K�ڣc���U�7�!�?B;��*���tvX��ې����W>��F�nN�ŠN��������ytx =�IM̀��"p����-�?h`��mJI8�1@�<9&����)�~�ظLǌY�$���3}�#Xq�Q����LU����,%�x��a�`ύ����:�s�z֬�k~E��p:��d*)�`�AM�i�xBm���
L�a*����~6��l� Sˇ���� 1{�M�Zj5���F#�+���*nulFw�ƛ�����H���� ��r��L󣏖I�kqm�w�7?���^�[��̡e
o����;LPLi�oG�@�ڛ���&���N����gR�vN�Z{.����� `�g����?�c�?���Y�Σ�jM�x��y���JD�fZQB�y?�9��B��F��S{��߮�����j0�J����dn�$o�W:�kw��"�B��Rq�&n�Ҙ�{��&JT�� ��|�CS��)*��H���._:h� *��5f���"@�\h�"��M����8|����˷b9r�v��+��"�:%��^�r����	�\�(�������,�t&���z �j7�r��$ڤ�b|L|�~�������LB!aN	�z]JPm�s�h��x�]m�S
��cG�W�ҳ��?�+��:�����&���8����R�4?ِ�uNqJ��~z�i�P[#O����n������v�ܦ@����.��Ô�4Y�����d��U�t�d���[�:*�Ѹ��v����Z��=մKDIj��+ZHi�˅^��
e��-7?8;;����U�Zw����cK�Er/�#��E���;<MF������k�<
4��ܕ�sC<E-����RL����K����F笧�4:^�zza>)��̏#�oɴ{�X̐ikj�b�����io}���ύ��Q��b����9�0����P���+7���t|+[rD9�64/�C׉oOlw�}_T�Rg,-[��p�9�<��g�d�+>�Ķ0�#��N�A��40��v�ދ���Y��F��s�S7�d���nߕe�Yƽ���}�d�)
ox[�6�o��c_7�3P`!�+����k�B�m|#�I�|����W��e���|� Z�S���Px�	�f�a�0����'��;��joD}�4LE�	i��Tf�p����hX�!������}�<��;�[2<�=q�I���e��x��Q���&�Y�U���Ȟ\ncd4����*�����^t��|����:`B��]Je���Z�$�*��/����ՆӁ�g�K��&�]]<���ˊ�--#\o;�7���&ja���u,�f'_��#�Ϯh����.x��������������L��,��tN���b}�iWN-`�lzB�n��~����E�j��b�P?�Ι��.��OW$y��!�^o��{ܵb+WY��K���V�5�� ��k�)Ka��΀���� j䕳'�C�zB�]�K[W�-�H���A��)�tXa�ȷ��N-d�%�J�ؑ���O�b�6'�@��D�U��	j*���v9�<�5.�	��K̐o�.����-�����Y3F;�CaYJ��o��e���;�&���7���>N�)�@�[�ע�ʜ�;�J�t�[��
�:d��>��{�I��>Ȯ�.[
Knۛ9����X�� �����ج���v�t�-T-_YĽ��Ut��~�fw<@���;
ø��
׿3�.7~�}~��u�7+�A��W�K�f���E��'evb�z���DF?Ye�_=��#a.��[4�a�;�3W;d9vO���k5&�NRNC�o@7�3�;��asj��������ڛ��~�����V*���I>�u��g��)��Ll�;�h�:��u��oY��z&RL���;�ø�ӆ�'5��4�NkL���h�0���gY{Rc�C=${�DK��p#�!	�޷8nb륄ֶ�_�FIZ���i��P��e�KG�.��j9B3��"�ګ�o�攴`n�2�P7�=Q�����Y��Ҡ2�n~��dwس�6�bY��3U�FX5>T��ǟ\H�m"��0_��CV�A�=Ƕv8�a틍'W�d�/�i��7�_�(I<r�6W2l�I{�yB�O��\�Ҫ<t�.]$m�9��~�J���Gz�C�H���F{IO��=��2P6^�ɤ�9�A0А�*�!-M
����޵��?� !�YI�{��f�U���p�ulJ�Tȶ�]N����x=G\�1[/.xK�ˢ�>y���NS0�%�)��O��c��r|d�������X�!�5�(���s��Kj����}�h=͠��[��5Z�+���w@D6���l���qHj,W�M�V���u�x&�/�x����~-0S���Kz-��T������N�����t5���&�j��W����2O^jp�w~�_�8�m"�t�Z��C����1r��^+�Z�VtaӸ�lԉ�Z۵�$��D��S����7HED���Im��<N��'M#��\�#]�U�|����	�:��e)�)Pp�M*A+�$G$�"��	}�~ja���2�d��
?������m�@1/O!�3�bҩG��a���b���R`�ֲQ1���%tDs�����Ki@�u�d�k�n�xQρ��`���a���0�Y�������a���t�}�x�1���ʌ�
��*�~��?�W/Ϣ�An>웮��g�D!.!H9aG��_6�`��
��,7<���z��i&�{�����zZ� ����ŉ�����Ҽ"D�.]�zc#yG<�,a��z�����x@�i9/�('��A���2h���a���Jɕ ��,��"�{��A��l���s�[tA�+BjǃY�pNԣ�0W�G�f�$�{����ߌ� �:,�4cC{�K&�lz.���%<��n�C+f��k)���:}Z�^8�:F�����CY�J�q���<S��w�����I����4E� �8#5&�Z����E�t$"E���P;=�q�<�� o���ă��3�
o����eAYg%?<O
'J�[J�3�n����
M�4˒����3U���O�,�iٙ���v�?]�B��}�c���Y�?�p�ԗ��UJ��6�`,�=kˊ��C�6j��e,�u���y[���ȣ�[֪d�w�cs_^'��eM����ia%��՚qpc�:͘��p����`W:�t#i�����@
j��h�u����C�F��(�{�֙�6��ɸz�|���B����a.I�j6J�_��|I~��U7�`��E���*p+�ퟠ��5���Y�RLzj���7�@��K=���ٳ0�qױ�4��X�
�B�������?0@+��J&�F�W��܂1�X�� "8�\.�Ʌ��>^R7af�̨�
����]��~����T��ـ��K�	���Uy���}��]�x�u&PS��FDVivZ �uJ�?���E_�� (�w�'4�03����|��,F}������L�rk��?�Z/���g|�S��2,���Y��=i��Xe�=��G����̯��-b�����"�g�/b�f�Ee��B6�g��#.K�(���B�lG�b��7�UV�,B��ܥ�Q���ݔt���=��7��������h��Ւ���ߋ�7@ �Q�}2� q3~��~���KB]U�q�?T:z��1�ao%�I"��TF���Ό{���	����s"��b�3%I������!F@mpbȾ3��Ikwt$I��W�������xz��}M���R7��S���B��l��@B�/�l������X�s$����4o��0����������0¸���ͨ���ER+�{j�����qL�1xѠ�|(c.�{�=���1~�G0VV��ɩ���FBT8�jޱ���>rt#�X�����c�=�Ҫ��,m�ԛ��OFA ys{-J�Z���r
(�Ek��~�l=I�Zi)��W|�H�b JbKN@ڶ���XsC�*܋ޫ�1�_��[���O�
�O�gLm�A�<UKc��h��l^���
�g]Ӕ����?�$�^s	U|NG��Z��>$�5�I�����5b4��������\b�d���$Lq0������.!Lk0|�lD�ѐp!Oc��K�~_�{D=M�L�����R) �����LR+�������<�{��0��kP�V��] &:^��umGC�3r������Ȟ��w��zb�E�4]��~ �?��a$���bG���+��.�yx/��WwE� �V�j�NW�=��9ߍ�W��o���۹ā:Yy�� };����jv����Yf��h���D�����n�bAC����٘�0B���F+��QD@�d�4��:�ykX� ����S�l�M]������m���}�H!e��̑�"Rd��c��#�vc��cCq��5�Qc!B���J��F�)��<���-�����~x��u�=���J�MM� P�{���[�G1��3$y�� �.����>�E��(_Y����v9���N \-� �$1�����7�L
k5uܺ�/���$"�Ne��F�=,7���3��I�d����R���#�߲n����p�g����l����Ѫ�C�Zl�(����ʞ)����~�;����E߫��|�n��t��Q�+���.kl���D�Թ��Rz����1���upYu	��X;@��إ9���nd�=�<�8&g���(���'�%�a�ҪbK���H@�����t���p��%左�za뾓��F�>X#,U>:1��,���&O:��C�*�Թ�i���������3g
[��p��.��8�k�������X^}dfl���R���<q,v�\-��@�(������������>�c�V�@�M�k��A ��#߷w㛾��Q4���+	uB�W��Dw����y��O������oc̥�p� e1�cU���2Kp®;bћ6��k�h��֎��Q&��s�D 8*���DMӖ�"�QC�ߠ6�Q7��o�1�� �F������Kq�G��GmrT���d�L>jY�GtTj|c��6�.�EP���^��0�b�U%���_�ƚ�iHY���x���� �� �4u��}�ʳ�\�Qp�s��'���#ٜ�>�;i���|��y�>��2������,��e.�ï(&��"�i��(����5v��u�����]��� �zc�u�o�nh��2�F55�ZҎ*���N$ꬷ����SҜ/|m1����I���~0W��9%/���������I���4�`�h���g/Ŕ��=zKP�f�Y��S�'&�6�:ab��Wll����N�2�ND�.4(I�ʳ�v-�NP��-�?���XS5���ǃ�6(��M�|�Q'�6��$�J�P�6�+cxk��Rh���w&���Bΰ�������/�~�#�'����&A����l�0M�CD����7^�,��1;����(%]J�dN��
	K���w��)n���%z�?��ŕ]����oxh�3�i3,���]�Ҵ��K%6B��<����82{d(b��j�qP�T�AF��N��VQN���'VJ��?=*D�$yyG�_�.�8v�2cQq �'n6��g�I�N0�}�q,�?Ʒw��1A��k�F�ly�@��ZG����jޢ��ڈ�?G��T��ΑeJ�O��=��M�L��?~�H��?@-��5�砕�L&�;�=�"F�dҋ�w�B&�%xG3ކ�NZ:�_9�Gif����;]$a
E���>��Y�(�*"���p?�Hy�԰�p߉dv�0b$@�_�ŕ��[���U$φ@6d�G$���ўN(��Ƥ7_i��
�;�t��(�[K�@c� �v+�"T�'k���C���E��	��o�ҥ�n�n���0����Q�]�k��~��2N*��y�-��Z�8�8�Ɲ��?�	I�im�����}����ߋ�tW���H���p1f�  �͋5���}�֍��[v�kKZ�7��&����ν+]���Ͼ��`2qJ��0��Q%w��ѐ��R���0b`����ͮMd'3��}���w­�CQpŀQ{|�k�:Z��;<����	�_}�~���Ƒ�4!���_f>3[(4�5��cb�3k�s�K_k�M�M\����'��F�2��%�,(��̛�TS؊6��^2��ꐅR�J�hW0!$�['��-+��E��{@J�>�����p�BY����|�9��a~tB��AR����입\�5�'Ի`�P���]\����8s$��ތ�����\�hkb�/��ͺ�3xRS�[A��\�	��gfV��?S
?��������O��(�9���{̜ɇ.q{0����Qw)s�:�g�	7F\4u��+���>ľ>f��)..j{Fn�"�Eu�c �����RB�)�D�v�R^A�r�D(�8����/�l8��<HRƭӋ�Q�N�����k}�����P�o+4H��r5��V09�}R�m�Ra����Bv�6� �pe��gGp��{��y{6|6f{;KI�R��>�.��Iw����Dg�T���a��(�i��e�Q�挲��/�3�7�do��.1�͎-P��wY���	��s.v�1/��	�׎����W�a�ũ{�{���{^�ںۯMzx��V|��f�-ݳ+D�?u���RӮF���?^��֯���z1��o�L�Wq�M��́��ף��9�d���\싶?I7J�ҭ�4O��6
���+��S�$�2���������3埭q���ߊI�ޞ�
ܢ|n�oT�Bm�6®]�����hZ^rw���#۴!�ȫ-�������)��+�p��:q;�&;��j�(�4�;�ţ��@���f�DH�����x�>�R�r2�$�~"�P����C0B�J�4�&vT�
>4B������:���G�y�FeQ��W2���(���%rqS�w6�;6��]Rէ�����Mh?L�j��6W�����P�Th����O|�C�2Fė�f��V���	�QV�����F�G�[�Jy��y[3��-Ȼ���?��N��r�e}a�Wsԍ���#hb3�� ��'����$o6/~6�/T�毹,lm�f�T�۽m��UG�����arI�9�I�ӑw��.��qф�ඓ@��o(tM䈨� �4KL�v	�7��	S�{���ܚ��y�A�OG�b�n�[��Mه�����0@����W��9��5��[EU'gn���,�o�'�eU��*��|oj�gr��������~MZ�YD8@���W�ǳ��Y
l��� `�u�"W0*2�6��2.��_Ǟ��yO~��������8�nV����n�i�L_��L:��␢��פ[1�����lu���wSwzx�}c��69P6��J%�L�8a��	z7 d��5�~'y�N%O6�'�p[P�:�*��B8�vL�6Yn-�I7�T�u�:Ex7[TL��\��Bo��
�t�JZ_8���j2�+>�9��$�J��Et�a2�$��@s���-���2�	v,��}PO���.5�̅�X�XR/��/g��VzYP�ye�-��}yl�.@��B�\[_��G�R�L5�{�<��[��i�<=���y�m�7�4�[�6�[s4 u�Ng���5�[�wDhmU5t�*�v���L��{�ee��]�ȷ3ȕ=g�ZD��_	���jx��p�d����"[?O�ܘ���O+�9���G���U�]������my�K��9������D�QFm��NxyC��,�rk����u_�Yw�q���n�U%@��7}l��_�Q���K�ں:��V�،n�u�ȡ�h���(˽{�d�4>��w�(��Y�ֳ7�.��Y���|.HUl��a��V�խdA�P�Sm��	����L�Q����
W�y�6|B��v�i+w���;v PD�������o�ڦ�����JH��P9��ͣ��@�ml2�w-EJ�'>�p��i�T��K���1/�9�!� R�� Vz��¨^��0d{{Ga��°�r&á@��w�x���}P@��P�����sRֈ�[k����U�ơ��>���2n����9ݪ���Y��P��|�{�����x �S�ɼ��&�-Y|#(���R��y�E�gM�j�)-��B�a�P�n��n��~,���u�!�*4WlwV�q�/���Q;iE�u@&ؽ�^��[!�q;W�+F����F�a��	����aB���$�Ӏ�㠅�Q�_����j��7@ 3 �nR9�������A��]���#�o�k��{����h?f���
���}���Ө�H�	��6��tZ^zZ�8�ۙ����Oe1T����c3������O
/�e��׵o9l�"i���n�י�gmX���"KȩqeS0G	-�ڔ��e"eou-P��%mӓ�Xk��=�0���f1��cVe+��3�y�n=�����?khMq��V��s�86�/}���T[����K��6��d��wa�wađA��n_�����#���Q_@:�7,`4��x����Y:.x5KO޺@���Q95|��;� <����ݾ�ys|b5��zD|`f�3+��	�(jN`^*>����!­>���8�6�"d�y1��i]���>;�ύ{�9GJ��*P����n��1+$U�@@�8��0����V�M�x����ހ�H�#:��c/DZ}Wq�y��� x/$��������U�����5L;���SA;��俅��$\;˿��*�b��$z��~0�F��f��B|�y�}cR&%��:� ����$���R�{�%���6���m��9�����q않�����KR����TC�>ݛ��1�մ��ʠ[e��.�z��
�L�ƛ���Mĸ��<���tkT�g��髉)�l���Z!�0�r4�u�L�
��Nn�3�Ye3�?~��.��vÌi��kz�
�p�YvL���9�U*lI�-2`T|�P�z,������۠��g�Ac���>����x�m�{�~��L-���<�c�K6��h�!0B���L"l٪��*�Ei�.nR��h�������������I�x�К���:���q/Gq-��/)�q��Ї�+�B�.�[H��#�1лP
�Me��QV)�\��d�
�a��8��[9y�{:k��͘R��<g��yb���K�^U�H����Z����y<��.�P��{f�o^��s�~|���u/�~�F3n�\�=���N!$��\u�Y���� �T��+�<G N[̃��C;q{����y��l���Ak�4����&ų��o���#䠎Y!&��.�Wޝ�
����isM-Ƃ�*��nN��u�3��s�V�G/��6�"vR��1�A]z|��g�m�oȼ�9��:nyC��EL���@�U��iR]\�8ؼ�~ ���b�Ɨd�Sy��_=�;37��v�'=��=k�U%E��)�De�~�,DLRh3�
��f��A��=]C�*��a�Q���rz�p�{�Z�p
Tz��[z��!�mmE"�r�&���ɸ#�l����p�$������ɬ���,���G+���?��76����1F;Q��9Lނ�xl7��{���xzn�8f��VFf�����X���U:p�Q�A��Ȍ���4�_#�y!� x�Dܮv�Ǩ�whR�
g#�V!�<�Em����a���m�I�Y����a.����v��aZ� ��)�I���q�%-h;e��Fj?)��5���+.��M�vu_����Ҡ������̞���X�a�AiX��ݝ�T} UV�7�a�Za��&���z �߹C��vi�԰����k�9��'���.mq}íct�)���VG�9x��Q*q3�l�]��jL J��G;GZ�	��f�����e��O�,�y���xO�+O�hx�ژ.;�[q�*����#rF��2%jf^a[D�w׺4Nw�W����\��Eeaa����y�U�{)��}��z���貳y���xs,�^�µ�����u&�(a��"D�W��-/��)��	$DZ�"[�|��i�����la�R&���o��
��VRX!�ҡ,��~��JM�N� d�j�<ލ���2v`��6-gp���L�5�y_ի����kn�!��V�]�n#w�G�k�Ľ��4�X"��O��(�]b�2�#;=��ǎ�b�a޸��!R�`�RM9��F�R�z+�»'����>3�}�4s}��+��ă���Ԭnnj�����&2`f?��dՂ;��v��sg�V�����6�}������%">G�\u��@N�V���]ڷ�ۮ���&�ʿxT��������.���@��gE��~�Nk6�ۉ���xUڹ!�~�w�(#*=�(�7մIEM�yk�~�V�B�)���ֈ)<��/ﺇ��1T?�@7[�����|x��@K��;�'i�&�a�nM�
_k�SO��4抩)8*k����g�nyp�3�4��.��4��9����BT�ۼ7zD
���D!`,���3Em ��+\�q��w%�d�&�m���*�/� ��PO�� �`���Ѓk�!L��=0�8zGV,�G�n�a���a'���D���5��*�zC:�^-9S�l_�ȿU1g+-�-/��܄4�Ȧ��Q)�&�7��
m7���������L4�0-�P���ޭ����� <6��a�d�C��v�n{�C�P�
�=4��N3{�m�4�H?��	�{tz����;�Ba]�(��W|� �4*p�� u^��]�Z�׎�/��¹�����7Ą���XŰݠh����_�N�� �`���Q�.��>�x1eT={SA��������\�U:@;�k2�	��,셧�	3����l��k�'��y�<��YNt����{� ���jNjɿ{E���=�얫�ʲ�9�n������Z�e��k"#��tE	�\ݎ�L�� ?�3����dk.��2�ħ�&�R�u�u�й�M��(��ƿk�E���<_�Ќ,��۷+e;��N6f�����S�yl[�99z<?<~һ��9��kN�0�rXr��f&�26���hŎ\;o�7F����!�A�p�O�I֧��=���6H�T̆���� ���:٬pכp~���o�RD�6�9�K���#$b���j}8q��Q��E�7��f{IE���*m�t��ǘ�V.��d��y���E�J����
����	}��O�&[/_v:��F�����n���)�&B�E�s��7��Y���:�`;�K/@�E3f�j8�8,��"�[\3�F�@=ke��@8����8v��d���"ȜOJb�Q���ٽ�N>]rA%:_t�����fx���$``�}a&B秘�	�A�����L�"�J)nYE���ws��tr9���o�H��Z����m��*b��ښz ��V���������L���Jr<;�ħvZ��S3�h��cox2���f����P��8[���HpD�9Ӿ�(�{�ҵ�=�&��Ēۄ���gq�s�Ө�|I�K�&G��$�����.Ѫ��ݟC� �A/Uu��fp}J���g��[���"c�%�baq[��w+���#��I���x����7��ª6�s���ޕ�Dě�c�J�*��n*�d8��>�p'�L�y��������F��Q�M	���
od�BNLֵp?j��Dy�����hjWt�̀�&���m�HLs����#MB� Q"��BL� 9"e\v���ջ�Ν�#�7M����=�V���qS¤��Й׶�����.۾��s��j�+�o��Ć����6vN�G��l�?���u|.k��PRQ��M@��Ae}��������E{q��K
����ƣ��&&�JJF?�z_Ś��
��߄չH������Ø��szF|^@�l�j��u�����yV�-ٿ"zs�Υw�C���JM�O��u�<da�r�}mj^P*z,���$��GQbM��r��76
��+�k���Cע9�拋G���r���&�>�b-t9��!�f' '�G����7z��:�V���jE�/!����=�5]�bc�3��l�VkeUpM��O-���+,[��$R2����R��v���*�[���ۯ
X���
�.bߍ�z�￧s�+"2�~�(❷�W����z��o��T�d�P���V8���\�V�N�$�n��8-J>Rn�i֮U_��)~7���cT����C�3
�0���X@ c�s���䆟b� �o;���h�s~�J�>�[x�e�La�i�c L]E�}�����{G5�u�Q��Y�-�H�#]:�j�)UzWB�	���M:��� ��J��[h�J�p���~�;�;�=㌓12�h��,Ϝ�y�z����MZ����,0�񠜖G.`ʡ鹽������}�g��g��"�LQ�
5-[��aF�Z��vp��q�uxz����;�B�2��5k٥͟2�o'�!����8D~n+�P'݀��5���c����_���O�N<6�35�hv21z鉔���ؒ��mN~���f�Q���!�4���vת7���c�O�!�ͽK
���ό���6�.k�(&IHxm����M���-(��S6&�����ՠ�v� ����,4I��
��0���qЭr[0���s�#F���q��ژE��L��Q4Pa�����b��g�&�>��[����,!�����'*��n@�K"�#�{�\�#E�Q�=l�B\���Q�U�ςK������C�lj*�L�.yk�����M�	����"ǻ�EK���A"7E3�bKNInmP��=dٓ�O�1����Ј$��Y�Q�l�	���[)$M�/����Z��g��vlzrV=͙J�i��x�,>��Q�F��E�|cRq�M�D����}d������X��o��Z����2��lR�b�gZ��b:�B�yD�������"�L\�b3�m���<dǺ|g�0�$�E5��2�&�S�?WT�=n�8BȖ���/	���XW�M�5�LQ�j������K��p�^�oI(a>��G$���D�7��Ǒ�V��4�4�	�H5f녌��:%�����	̹�Ug�6�A��y�h���򥫶�\F���8��ښ�Ι�/ݣeӆ��@ꂶ&�,�4��v�=�c��s�؋�Tvםb	�}�S�2IB¡�o�O��2*mQ���3ffajT�"�{��)�	�8��̕�꧉z'/����	�b���t���t���L]|*��d����-e��˖� Ex�&ս���nؿ#���x��BC޾O�k	��ur�����l�x3Y� �Q+lbiawD���`��(�T_�M�s!U���͘/4���Y��fh�Q�J�&X����~�0/�?X�����O?������y��	� 8���ʽJ���1�ܬ9��G(�XZ���I_P�7%�*jjr��l-?�7�����W�O�Lѭ'��k��YaL;	�����ڮd���O����h�0����Asa9������?�2�����w��":Q�b�Fb���G��tT]�/xl�!�����s��O*�Fx�����~�c͖���)����Cc���k/щl�H$~��ô����ҋR�Ts|>�N�_@��ii:�=�J��/Gس;�o,��z�+I�SL ����c3�.�t�]�k�>KE�
!BCo�Ѡ����	*����%I9�?Fi+]uǕ�.
���qf�������ڸK�� 5B���u�Ĥ�	ӇqO�.��퇊<W�'�|�^!��g��75mthB�:�����਼����#��B�˵k�W�ʖ��F�Ћ�R�F��[N�����,�
��Yh$,�s�^�P���3��:7�zW?�싡r.�i;������:�|�;�h��FPk���A����|�;�����2;�u�Ȱ����C����ܳ"t�ֺ����C�:)�m(ܼ6��9��Ĵǧz���<>fl������:$U�I��Vb��4g���%���p3S4_;�8PN��X���g_&�6S��lc��X���C{{�{�}	�E�x���Y-)�4|�'��0S`�
��K���xH�<�%Or��s8�� 7�[��tX��bT`1"������-�l��*Vܹ�DZ�=z<Gu��(s�Z�4{�甯iG#��|#a��8ޣțGE8���9��L>�g h�����?EG]���7�_f;�L���u��pN��oG�������Z�o��B�EW�fT�nj�K+��vJ�:��/#3E����)	���	�&��o�����<WL�7��r�t���M�=�(m�W���������kU�`�ѕ{m�Y?�[y�Ŝ�Z�[}��F������V#��ֺƈ�z��gOY�`6����BPnO�L��3�^���Dp)V�93vY�}�>.����@@���jȭ�-�hV�A�2,�Ň��=���O�����=d��7�pD49�5��~�S����������斳]#�b��\KNV�u��HC,g����T��6U#]�%*�ʹ��^��!�D'*qg�NТ$�D����z/�!�c���[�OzD�
���^-ұ^��w��,�v(�@;|�yY`kՉ�������6fX�v��$�λuI�.;=mނ�9T�ѣЖb�D��=�[Ȃ�6g����q>Ŋ�(ӫ
�hf�ց��DQ�Ѱ�{{o<��9���=���f~*n�D�C}������h���9NI�����$�##qUȄ��;�)q���h�A`|�/]���V�� �+"�Z�1»g<�7+0�u*1�7�����<�ˍ��ա{�=Eb�[�����Ң���.O���l� �*L���:������V���"3�+�~t�k4�#23s���� ��_��������耒� ��c��`W�,�H8��2�x��!st4�+So�+~�<��#�py](�����(K�5��NK&)�.��9l�Q9�8��O�73#�T�^���*2�*+w�Y�Jt^<+�xF���kdx\�wn��c�u��{C7���cV����)�!I���XE�|Q
<[����EKs*���������Th��U���q��NB"s��2��P�퐽�Z7Dn��	�v?���*�~���X�^��R�7�"��A:P2`�=w�?cwy)�A�PMucfT������)'�gN��\�ϝx���m��ls�u�H�u^�`L�V3�'���r�)�CF�?x>�Jl�"�z���Ō>�4��ZWc܏4,%f�������~���ѷǗ֯!�L7`�z�#�u���o�!�$�?ʴ@��(_��y�\+����L�#�V�oGC�/ߝ�$%P�����ld:m�ҊeF�:[W��J�I[cC�;!߿�d���7��z�%#4�u��s]n�zS�)%�����!��d��r��Us�@&_�EO��~l J�a�pd.��:F���y������&�.��	(���i#��Ԝ�$n�����=����[�����P�1�L�PX,u�O�V2�H�%��.+o�1����\�B�Zw��Jt����L��B��F���ƚQ�aX*�d���_k�M\�M>Tڴ�"4��:�mP�c�����_.]�\eQ������A�ts�&�o�d;jLga9	�\��>�b9��Lֶ4�Jg'O�W�<P���8(S�K��d�H;vʡJ1�� �yؤ=�r�˕$�Ŀ����0�G��>VW5*��ۗIB�r㸱�K97�?�&:����^ Ħ�h��o����7�E۳Lk���͎��#� ��T�W�[y�y}�j[|$�4���;m[�����N�)��b��"��*_�6W�qf��&�N�<�^������; ��XND�@��tK�����Eq���?Ǥj�Ǐdx���N��a����kU�.f&���:�Y��.�6~@���PF7�/'M��G?iX�s��%h���*�n#�(19��wX�B,�0����J쭂��AM�[�i��Bȝ�99�0���)�CGQ�h����G�Sj�T̼Q�0ÉW��w]���Ff��F^E���~�R�V+σ�G���葃ھ��|@DW����Ն�k���/銶���,�´��Ŝ��/Id?4R'��pn��o�]����s[&&c����&t�����T��sv,)�:�:ĳ�q�'�[�'���4U�����0��g-����sҾdf�[AG���g��]�̍{�ڦ����c9-�M��\]jrM�3�z`=p����_z�8��B�ɳ�h�+�\���G@��+X8ZM&�����:@��<��(�m�x�_�������$vG�:X��$�y(�4���2%����]�j6QȺ�c����9�3'%��t���@s���jF�ӵ���o�iB}�F�����u�U����j�md08#	#�Ԍ����t��%gE�D�rx�9i%�(��[՟*=���V��n�}�\��5GB�:����J0SG����gp���!ƀ�'��
�����A��yc��ŋ���DI��$v���4�c:�Sԫ�}}�W���a��0�������.tO��V���pn!�w�κ�FQ��"6��$�KY!�ysl����_���r1^�[K4M�0�6�-������x����c/�Y�ùɬ�6����e2R'������9mJ�ݷ�QTMN�=����}�ﴷ�Ѩymڂ�_�=[�Xx������w��y�"%?��b�T�P9�I�q@J�V�uGJ���X���^����yOz1I��>.,�=l��:F��K/�s���7�m�#"�����1��ߗb_ M<�L_V�G��*�ε�̡��}���ɐ���W�u���n`�F�/?�,�1�3����13���511�����ǐ8^�J�([O���ٷ埵�5��t8fe~%�j���!i�S~Oy��]g��W�V�(�d*��S��$�(w����m�x�5�P�a�O
��J��k���R�8XnX��6$hpD�m%+P��T�u������2c�4L�zVV�c���8\}�����w!�UO�кy�RjVê#��4��b� �2L�C'��tZoU������śƻ���Ֆ9����E��ME�w�d��S��K��#e,c��ɷ|W�Я�=�W�?,j.n�o!�@.��%.�{����!���͐�x5�:V�W��[%nCŅ��:�q>sQ���Z�8�y|]�x]e��=�m:�)I��:�n������RTj�v��m��F�^�����"�9���h�/�M�3�jR���4a�lw��8kt�5�86C��#���[��V|��?�2�ݜ��P���)�mЋ��S��Nq�|��r�GnYn�2�W��i��U����$F��#�y�i�OOO�d���[k�����k��fq�nf3t��S��H�B0#�|��	�0�~�F�8��N�>y&�̓�*���r$k��F)���
H����y����u�o�\�Մb�Q�l����ߘ��������V������� $Fg�<\�-m�| �Q`KnۙG�ai�)�?�u�z�,eec��zc�"��D.zUs@�5��h�5���c�mq]%��P��|��d�#�:3N�9�\��g�J#G���u���@G�x�B4�as�bV�����
ɬ�Q/��Ԣ_/�[�%���ɖ����2�zJ �j����\u���\��Ź��i�+q%�:�%�Y���?�:̜q%o|o�ƺik~&3�K�,��|��㬗niW�躱�g�����X�T��w��T3���� (�:��j���������p�歕%�)���x����EU�؀oߍ�r+���}~��|���58�&��*�#�r��ߐ\(
96�7Z�9Z��3s�� �`5��[��+��k���n�ےf�G�Ȟ��ėS�
���DUFE�NɌk��^�^x���?�;�H �U"pխ|������,�J���7J�5˰����;0ڟ�;=�"I�W�# �;�ż�bۂc�HCVO����y�z�����y�5N�H�!j2��o�^��(�-3�M$��ғ�����b��+�v�h��n����u��֣���N�|�2m�t�g�Q`e���]�b����H�g�Z9Y����!Y��XֹM�o�iЭ�TP펯�_l`��
��l�l+B��q~���ىOR�mH3�RZW�WU�W���x�r+���+�#�Ϭ�nq�}���P�rUx���}�Z��Y��Ӿ���*��;�@�1�繢x&]��uO7��7���fu����"�����l��Ap��9ށP��X��+|��n��40;a�ף!�=~������/Q_1_���B���5ҋl����}��6׵�oJ��)w��l���g��Ew�(���Q�D~������T�y��5,����C�cI�;E��]C|����sf�'���Y��3��0�y�(1��HN��s/���.٨���S�w�P�Gn�\��yge�;�!Z�=C�$q������X��o�M�����GXֆ����GY�󜄃P�Bq�*N�D�sؐ�_Z�~��GQt�Ⱥ��o	r�0�:�
�qr{;G�j*o�Fd��m��_��]v6�0c(�{�.�bضV�b�ڬ6�9��~3��m��.p`��������W��9�y=ƚ�E�_O��6��+h�^�`�8�c��%���k���uc9X1��a���5K�΁r��`�����hϗ�6�_=!�1y�G֊Y��a� PW߅)g��~�_����e]��7q>��=Օ%���v�`kQ�Z�1-���-�}VQ�kn}Ͳ�)/�e-T�̈�U��p� Wd\l)���	�Q=�j�;�p��1݌�>�Ǖ�~��v��w�{�����y��q�9�6u�21���+\˼W�EW���{Q?&�q�ZY� C���zp����Ĥ؈d�O�yψF�u�g�U�=�a-A���#�ޢw���q4�j]�"��Z�����zm!^�U�V�e�н���X�7LI5v!g�yl�eԙ��ۂ�2��75�rl{�q�Y^�l�;��A����x*���*4����.�}�^��,::�nw�ӰԃU淪"���J?rUrR�Z�A�<�� 1��Dα�D}4	�(e��L��z�u����cs�0��-.�lDu��:��w�W
��Z4��T�� U�k����xs''Pf������gX�$��]D�<�K���Vl�P_,@�mK���\�0Z��#{ �Cd�9l���S�g>�e�9�X�C�Y�6@��nYd�"�2��NO9R��o�쬿f��%�^A�sت.�A��/��m�MU�uu/=�y��tku��PRPi%YJY\���_�ȷ�![Ȥ/6�8}Je8T�@o�`�*�'�q����|3"�j�-`���Z�j�]�2Qw��nǲ���+ Zv�g���@� �ur ��IX���C�F��x��M2qT?���`��S�F�!��r�����jҾ)Z�뜏+�kv'�D�!Fٗ�ڗ#xM q��%ܐVQ��O%����K05h揊a��PQ��߉�T��{͸��NL{�MM$K��pZ�zc�Fϖ��@�uYATŵ���>H�%:�Ȯ��ch�_�0I`���յ�I��mF]�q�!�d���R��iM�.J����(5����{�m�E%�{W�����w�L �E��vs��N�ߦ��l{q��o`9kӰ�eN�<G�_����G���� ���Gc�aIq�S���UaSP��q�h���L�
��Q[k� �?,)/�������&K��t �� ��y"�|��@_B��uu{T���4H0�i�9,�<W��w�_������� �9[\��bDt��o ��_j7��{�*�1d��X��oXx/�k�t��'6z���s���ck�[����@��,��a�J�AMTFw'ݬ�O�'���9k5�c�*�05�|��H(U�	!�,�o�ھ���_���E�
�+Nk?�p���b��HT�M���*��~ -_@�U�A0���O?�mc���ڐ����:�0���A���#}FW ��3B��6���refAR�:]��L�4N�{�m��NՔ�S���=������x��dz�!n�����5tg}�!���b/Xf��*�l�]�!b�����s�كq����\ܒ7���GB�5��x�Q���S_������-/���@|P�f4*�m
��)��j�k7��h� ����Nͩ/wR+	�F�a����~M�_�V���� �>�,-��l�Sk���;��HY��ܳxڃ��]"�����+�mv_���U�T"�� ��y.֚zh�	���z�mzj�a ����&����Y�k�xQA������Y�Y����A�W�\a����� ��dr�4���zU�bNe�˧�M�>�+�`�vzU�PJ� ���z��pl���& �y�Cj�BZ}^���:s q�:��Ζ��蛄�h�q�RЗ^�	G�i�Olr�Ag��i�}��@u����V��7�� �+�so��7c�Ά����Ɩ[7�sFs�󹦭�-7eH����K�;u�i���Ǯ5��/\�����m=�#�A��@�L�[���A?9H~���J�v����)�*5�3������*�=f�qEbq�t����N�p+KH������:»�i��������3�6��Ⱦ7{V�?���B"���Mt2[A&��J�Qm�_z���EY�e7٤��#���\B��:&o���-Ӟ�K0��4��	����|a����n�t��=�܀�
|��^��9���Z��Ux[�^Er����m���I�.�����A^ ܎B浟\Z�&���a���EO?���z\Q@��t�/+:�'�i�cQOa[;�ޟU�g�r:	���@������>�!�ϔ�����҄�q�ޙNR,�eVDV��~�|_�Z��ԲUR�z�v���M�uD�&h0Q�z��u��h����<t� ���	�|9<]u�;]ޠ��e)�d@_-sr��w����T1�t�V����e"=��/�U7�{!�% �d����y��P�A��?��.�ʟO4����ȳ�v��O\ʭJ�b�$Y�b��#�޸�`�+��]|�@O:Yؽ{+���x%�b�ͯ�
,��Q;�Y6�?Ы+ˬ'+�Va�wԋB��O�����r��(C��>���&hJ�ben��'�s?~�`���K�l�mvO�vz����]"�[����'���>y ������p� �y�B�����`�G�!zUJ�o�i��$�Mܣ��`���poOF���M��Vc��4RCrC�5�Cr��4�8����8?�ǘiվߵ��*����?.���:�`��F|C�wo�>|�(��ߺ�S���b��U>Q������5��-���;��3LI��;)��7k��v�R$��dM��"j���f��VT�V��Sy��lH��ҽ��S��oiI+��p��rE5�+�XN��Z�������x~IOS�l����J�tI�鲽�~�Go�&) �W�zm�^�<ր�����Q��-�E~spZU�@T���Ȏ!3�}�Jc�H*�<o��T�2+4(�����aJ�������&��V��:C�+�����U���oA��� ���e�.#���g�zf6��U}_�0�3$p`���{�st�`�؋�?0w����a����-�ϏO�jd�E���|�����]�lX�Չ�Il��G�ɗh+I@P�-q��9��NTO�a�Ǉ��O/���Ԉ82����霵GZ���A�`[��N�?��e6N�T���)Q:�r��C/!��bN+햆���g��h��0��[��:���S���/~M
��H;��}1vw�sv�:���ry����%���2����^��u�|0¨�nS��J}�#��<�
>�}����q΄h�@�GdP%x/J����{��b�[�9��~�b�FPr<���-��|#O�㓔<���y�`n�}�O-~3��NL�Q��Y�^�( W[#�t�A뾆t'�����kQ��Ne������w��#-� ;ˡ����l��������)Ub�KH=�a�-7�jѠ0���VP}��L�ʉ��7�0P7Zi��g�8���p�����E#��1������w��qC���Y�Lw�|d���B`+���t�X��vO�j���w�����EL�J*1�
�C�3\o�8�qX�V��*��(1��D�f����(�g4�B����I�����G��T(5��.A��/�yK1�l7��X�o��`F#1+�岺y2:zb�ͭ�iC
]�'�����8��솧��k^f�b�_���/��vm���7>>�:Lg@�L'����C�dkF������7���e�>�'�3�"
��X���A<5�&�����d�� ��?�=P���"��Ff�?jw�I1���ub���� ���n��Y��ҍ�H�4�x1O���]�Y�N���D��~�\�<|j�ܿH�ߓD 0���~��y-z�G�_���O��SW�R�^���m����'�>�ˈ^�9:�k����ubQ��w���۩f�)�R��p�[߀��t	�hNY��?�{��AXn�5��,��o��
QJM'�R.��Q�<a���}�X����7�s��>L�����~����[nO�0���w��m��U��E�//b�I7-S�HRˋ�-�-�p�'Ol,l���������7�j�?Z8.���*?+tb�O�?ƪ�(��UՉ*��z"kn�(�-X��z���J�b�����`9#�r�bW�H-O�{~�y���4��ZC����*Wdåu�z�LЅ�6068�J�g(�.�cz�k��Bxcrq�B�����^�}hP�N�K�����G�9J\��Xa׵�n��|}�!����W���!_s�Q��<���1�5e����&^�A2��J�� �K[�8�hl���1�0�W��	��F�j�p3�V� �k�0��n�D� ��8���<�Q�uG;�H���B�wm���P��w]��箿���kV�wkӊi���}�����mp�V����_/=�17���i���et��\�w2�{�XXίy�d���H���\[�R��wɼ��{+�<֖����\jj�{}�k�c�*6��=�Q���!>�@�Q�L%�`>�3�ݥb݋��d��y�ӟ��A���ug��P�wSʀ|��y�sN�	����i�0��Еc�u�(�j��k��|�\�ht����T{8(m�Ԕ�p���v�Z҂@��������G�h�s�Ӣ���Ǐss���3�������Y�܌sv�d���S�q.�a���TTjn'�V���)U*���a������4b�R�%5��;�up����w����z�"$kl��`o�-q�Z�Be�_k��m�<V*�ZW��0u7�����P@9�T<�Q��v��7�ǘ̕��7,G/}��gvWj�>Xޙ�5�3��7�{zp��t���罿77�||�|����ء�0��F#���E��5
ލ�2�ܣ��_1{_��qrQ���S_Ť,�_��ݟ�j2�(�o0���鬠�~w}�a<%Zo��s�qk���.��==������4�E�pr�|"]I������C��� �+��Y�j|9��
�L���^�}���O(*qP���Y}+suR�R���G��Ix���,t�o��C[�����0���W����Q������yY;n�9��h��� ��DG������}, З{���$Ew��8�R@��=$�
)�������IGO��I�߶:�\n{�{A���^��bt]R��$:9^��R�ҵd6��x�Ƌ�Ea����n6\�~m;a� �0����=q��)fp!�r�ӥ�_��q|�r>oa��MGl%��ٹ�@�j��J��!�}P~,[X�D��5�-e�dY��Yz�h��J$��n�o#.���A���DU��8Txy/ 5� ����n2�lZk�!���yC�}]G����N���͔�y�ڎō�T��/�c��3\�"
��V�=Y �:c�#x��������؎eoG�ݙ������_����zme��Ѵ�Ԩ����d�����@Gg@8�:N��ᶝ�0�w���E���}!r�%� ?�L`�`��_���v����:Y}w/c��@��tB�L<���	��)9۹�U�|�N�+s0���24b�:ܭ;tJn����=(��y��Eq��l6�N�yYyE}S5�l�c�LKO����{U#�ijU-*0q��&��L	�g���(�,� �	J����ӌ��,C��WM;��
��?�%�M���o��P���F$��-ぽ�վ5�����	ST�x���'x��J������c�݃�)���
�ϗ���)ɴ�u_9z��-�]�М\�+�E���Q0���nB3[�4����`�������f�����kv^q�T߲g��>���2�����j�=���Q���`~-�2�؄�=�n�11N��
7,k6?qn�/"��N�3�����p��`�K4�^qE�q�v2�68�9���t0�l`�����x�쓼�M�g�rF�4����� q2_2dPF��w�~�ʬ܏��/k1�=q�|����������8W�j�K�U�h��a`ŋA���y���S����x�r㶗���O[��8��}�_�ǿ��df�7M��qQ����
��&����"*���@u�H�(�O�XGu�����C=��p�}�V^ۭ �e.��4tI5�CXl]����f�/kq���{-n�*7��L{(i�J'�L7�	�����/u��C�y�#�ŭ>|l��n�Y�ڥ�w��2�'1WK�4Al79�i�Ѐv�zF���?�ɵVx���4x�y���)y?����y�X�.�c7�o���;9a�[Ub�~���Ep��Z0��K�D6cP�J�V� )eb7Kr���\�˾��_�?5K�&���3���#[���b'���#���&���y�&>���u`z�IJ�Z�����9Dc��v�(V���C�0�^�닌��%���TA�O����H(o�#��=��\��% &uW� �v�Ϳ�A��{()�|A�7��u2�ݾ���Q�9F<����jxȏ���_q��|�·�����΀:�l,�5�ޮ�.�_MZ:!#?�ċ\���Də���qC�d���d��bH�J�^�1������bO�#�h�:��I��G�sͺCC�4G7�=aHk��+'����c�p]�!�aM����.��-%�j��^9$5E�zY_��q�݅7kx�ᦫ�I�Ut�T�G����&����3��V�c9�O��U�*��.�/�ŷ:�?�w �ц�b˸�3�A�\2�/#N����Kf�u�<Y�1g�O��f���,HE�����+&_8��m7ڵ뫊k1�Pz����ĬKzl��MN�/qjI��{��6���s5C�(XfZ����~Ҭkra���['�iN�����ŏ�kza�&�; �E��Jς�?��V�!zX��o��)��|��k39G��lY���b�[�&N[[�^�ʈ�����x���[2������d;�.Ӑ�ӭ������i�����Q*%�жt��G���2
��}U�k��΍�T��r�k�]�by�ɞq�>f�H�~���W܉���O@�R蹨%2M>��41H�Ө=Fb>L��x$R��Bf*��V�������9�Wq��$�5����DDPF2��$�����P-�3�71e�P�^!�H�����ݣ����o�mmgdT�Ϲ�t�E`� �&m���H���@[$�л�K&���5����_�g�o����S��6����\1���8��⑲l8X��k����4J��8�h��@g�� �V���&M1�hqRPZ<Vv�)w7��+��ig��sҴ��'
��0�H����C����~���D�ϡW^�1W� 4�B��k$��,��U�q�3?9J�:�>��υs�|���?��HN�
5��f���B���*�!c�("����C;	aJ��zZ���l�3�(lCcgk��캛
�	��+Z�.�K��3���SUWě!��pQ���s	*婝�_@rЙ����OC�?vĄ S>�<���kx&b��P�ƥ���u�`}�?��Q�b���	K��Q����/)�_�� �.u��2x��뵲}�Q���,aq���y)��C@�fy_��o�?Y��1��ɄTq�q� L����(�\^}��������s�k����Y�;�\�ѻ�629�Y�3L�?�l;m���ͽ1�;pE��Q���E��-[������c��=���v0{ZU,#���rP���ҟzu�ֿxM�+�p�}��?�R�}�#6�l$H>��;��}�\;��O�&�[Ȭ�9̸I��DÅ��>v���=�		P6F�E�'	�7���A�yǵ�e�]�,]h8��c��լ=[�q������傳U7�'��-�>�h�=]�RۺLү�Qh���n��J �����������l�(sIT;����N�q�q>}��>��7H@���{�%���"s��$�{	�w0�+~�p۹�� �MT���y�)Z�Iۚ�z44�������%J�u��Q>�j�y�+4cN�P��L�I^3�,�ad���L��z:k'�Ή[;
ۧ/�aGf�eϡ�A�]�k��@�Z�!c"�o}<\��bI����+�b|p�Ch�ұ
��v��J��AZb����"���#(}mE�z��r�6���[[wM��`��@�2�)%������������]��S�bL�P�X�M	\���̅9z�q7���lܠ�d6�'������q��������2O."�]Iv�ÖJp�fc^�5,�`����������A�R�zE/j��S�X*�:82n�߰�����ĺ��¶�ǩbQMP
�QW>L-��W���o:�OD-`<e��i�}[Υ� �\vb�k��enk$Z+�y$��R�FJ�WW�ǻ�=�C����q6'v���������f$�䉯����iU���u�齫���O�W�������l"u�4�߈ �ڈg��$�I���;�+����(q/J1B9��,[Sk���*���/Z�T�	 "�@Cy��1��g܍S!@�˾M<�#��V�N�0���K珕��͝���Z?4�h�������=h�:����B�<��;gQ�HO#l8B�h���f��3��GVf��4P]~�m�4��a�o��[!�5,�;�ʐ�yS�Q�5��H�<�}�!RC@�4#Eԓ�l��jab�u�����a�+]�}QD��ڝ� N����u��3��:L>�����X��hH�7&��{�=	��{�z���k�r6�l{]eN��w'g�r� �����DlRLT����7ʫ�+�K� �����N�?��5�3]�{>��z>(��(�(����k(�_gf'`e�ei�	�V��I�N������ބ�@�����ce���eN�#��~^��k�P,��}���� �ǽ���K'�"Y��u&
Cd}�w�iP�ڕn�)졟�5D��tׁ�:��0��|lQ���\.Ɂ��q�WX�h��	�+~E�?�XR�.{�g-V+K��q�QL��`����ꛤ=�A)d$� qȡ��" 0=��?��������m0��xSGR�$z�����[�Lp�kw���ӗ:ݡ���n;�;G����K����N��%��~#����v���91��x�5+���7�^�s�e�<^�M���%�$Nx�g����<*��~�^EAtep���($>�Ȁ)��T)��\��a+��!��^/�W`j�1���g!?z�%����^Wn5�x�L�|L2�����G���n���ݒ�yY�Ha�R��q��u<��a̕�5#�~'�6�_u��t_ԯB'[�Jf���h4>6`�?�x-�g��w�Z��Ш6��
������f��vIsH�V�N�F#�ɺ#Ėk_jX��/0����z����f4���g|�!��g+�'-�a�vE��3�T��c�J�+F������RPpÎ�ǆzk�':���˿����GQ��-t=i�����.?�8����&R�a"�*�e�_�s{��w�(�]E�[_ߞ�g����5�v>l�-z�[�cޠ��o(��˧Y!������(�6=гX1�����x�0\"�Sg[k,����CRM���������I����(4`gË�n�����5]�1�V�����gJ2Q�=��#��]��K�^�`�  Ɵ�N�n������Dؖ��D�Z��;�,��kA�gY���iŘv��;Ǧ���s}�V���nw���Ѝx�y����Z�h�c��o�M� 1YrU8�/��E>9�(��s󝸹=n�hNh`�uT�K��e�Z�Ybc�˪�C�;��8��9&T3��+g���!<T�6�j���JN�	Hx=�#����o �n'	7Q̚ݱT���$-w��^����mg��K��OT��%k8��aJst�5ϑ�ԲZά@q����Y�2?U��[�8���4 ��z�3�p��Ah䡞�{
;4
ޯ��*C��k���4����c�]Z��X_E����;pE㵡������:�������?�#�ѯ�J��w:��#C������#E���42�(p`�����j5���^��B�vxw,!�|4.f��R�޿�o�&���O�&[��3ʢh˩S��@��m����a��~^��fD��գ��rݭ������/*���OR��+����2Pmb��"��"B~H{��bm$���h���fJش�Z�RL&���p��6�S�?)^n?9��Vz�n�hWdZz�- &�e��2s�-B�TDa�ReYA�x���B6�|%��������YE��jk��O�����$�`~\��4�b���`	�R�A��ڕV�}�77�,�k��`R�Ϯ�q�a��0�%(d_�w��s�1��`�$E����qnt��I���Kq��u�#Զд��Ud�����zK\�}�"�Y3V�hOE����.��̆�+4������=n�m�zr��$y�"�D�a�9w������;i~� t�����ΏM�u�_jEu���5��-��,�F���eSU�$���[	Eiׄ���-GkU�{`�v��B%Q5�Yu
d�(����B[[����w��I#T��b��C-,K�00;��&��:��R}��[���#�v$ �,���`ђ�E�n�jԲ�=lY�ٸ/vv�6
�a��cg��r�ֻ��O�FE�K�~]��,oWK/x����6�:�(���͈�m#]�2cj�^����.Zo�pAੌ�)2F�mÍ�-x�� �vi/�l縛l/����C�W@5��������R�!!*�J
#��H�(!��J���Q" �G�!���L��ϣ���9���x��]�~v��?�������\��Tj鈨�g���1�s�4!�$��Tɪ1z�.��NL2���N�*=o�`��N^����W��z�\����k��uꜩ�����[�nk����M�d�p��7��@��"6�PI����N{|�u��\��	NG!ӆ4�߇4���y:eb��q���r�8fڻ�%��|�x`@cK��n����KX�7M�T�AD�,��P��	�0�N��Lq�`
0�$�Δ�gԹ��y���Ip0&��b������y=麤�T�>ǙB�;��5wd�׺�b����)7�˶ۛ�m��	ƣ�����^t�m�`L� �v<ꭺ�s��}]���3�����bD:��[�S]�ܵO�)Hѵ������{B��H����B��}#]�fiB/�%'K��}��D���M�s�����ࣳ�L�l=��� �=���(�:7�Z�����>#}OPdx��.GO�&��"���W/@'\����4'` �b��Jms#S�
[i���4��HM׾�K�:�<%�YYƶ��K��ii��<iPa�a7W3(�@�ƴ��0�s�h��"��5ϜA��8͡=66Ei�w��Xq&<~,m��G4�9��cV`�)[��ޜ&�3��Ѡ��BQ�d͡�|n�b�B5,��[F���ш���eە�yh'-���}(�4f=l{��!�R�[m��a��ic��J-㽕�`��R�f^�31~d|�)��ו�"Phc��}�����Փԭ�JΕp�7v�8ڻخ�t��5Ui�=�i<<��ڹK3^��l��� �v �Zvf1��5��y��T��&h�?����FY�EͫVc�S��ce����M�݉jme�%�q��^o6�o�,0�B��M*��i����o�yzw�`�̊�����B�]�gV	��D�g;�w	NL�'�V>�_bj��xa�����jB%D��&�����V�@'`��F]WHtLӓD����{��/�=\I�]��_��X��i�Eii[*��m͍����o%r뱧�R�'W��|n��d�A���J��&�>��-e���hr�=�[g\=��!Ot�њ@���D.[+���

�=�A��|�������J��AQp5+]�{�l�����c)�h��(9|�tY�J	\fڍ��C�p;�.6�Ą�?�fK`���5�3���{FOG'�:�hm�K�,))t�k���u�s�=H���ۄ�#/|בn4��۶6����8��V�^����L%e��o�T���Kno1,�����6�uE�g6�w,3�\b麌�k3�&��{����m�Z��F�͑���ϥ����S�2�˚P>>��&f�8I���I���B�)��k��f}��Y>#*
��e��a�;�{4xyEƝ��}�C���zQ�y�4H����aa^�j��Z:#����U$���N��{��n�YFD9�W;_�v��ڟ8u�U�f\E-�?/&r�-�z�~B�[~����AW�VZ?,-v=@�õ����s����{0���Qf.�;��t�k��`h��v��<��Q���*�>�,��G$�U����f�>y
�m��H��S�z����<e����u�
�� ��5�C�tf0��z�IX����g?=�bX�39@��zl.�+f�x���$gp._i�iUrɀ�`�2u�'�1�	��H�A�>�>q k�xw��?\�^�΍�����D���i�5T:��#+���E��,�z��o�7�Э�47��+=�Y���N�.�ۧ#�U�^�U���VL�*�K>J�g.�%���Bġ�#���٭����A�ū��D��v{8�Ҹ��r;�zPjmP�7DL��rKtV�_#߂g#sl��C� T��n��d�����F�S�$�A�	�fܢ�-��p�uZe�]�{�k���Y����z@�X��鳣�%�)!?�3\�dBǩ�#��uX&*$L绰��fG^L��)>�|�i_�
�1���h��T���I���b�ݶ�
�
J,�	Qf���}mX6��U����6i���̢X#ޞ6�m"M��eI�?��%8�M��O>�s�?�����,䲴�(�����|�m���o�
+��#d�elg�+���O�ܥ�
R�_l�SŌ�J\=�BYgF�q���p��������:�/����m;E���([l���$se��� ���xN��)O�R�SO�"���2u�;7d= �>*/�N�5dKܽ7�٣ڗ�+"k�}F���9�c������T|_����E���[hH�iAd���YT�
���-�<�V��cޅ�aߚ��P���{g������Ω��y;Z������A;FtJ�����M��CQ@j��(A��ׇ�e��Z���]bhpX����>[@�ؠ�E**�6^g�lĵJ	��5B	�.�o�\�Y�n)y����a���\t߆&��pjx�ﾰ)�ҹ����<�:˙��J�ܨVu>u� a?T��kk\&1����
��姑g����]_�@H�SlGtun��h��9�5F[����c�@{V�g�%��r�����=�O�{ڲ�!���MǙ�u���E��5�3:�]Z�5H�$ҏtҟ�r5kO[6�tKuK�:\4Kj\�ԩ�.����C�.�:ń	ϧ2z�fAM���E^�.�(��O�}8�9�������S�L�2(�#ص���O��s���Z�AJ\3vI�)2��H�2�sPb�/dB`��9UX�s��O�n�N_����E����dw�w�N4��ҹ�4�R���:�H�����e.�3�k�vԇ��ڱ?L�Z�@jp�F�0�A94��U�V�"`S��5T�\D���:-�08���f�#S���~K���#���u��o�,硢�V1�o�4iL X�Ta��}u�r�a̡F�کZ�J��a�γ��I d�И��o\gLl�����9揎�t~�Gn�>Ѡ5�>��Jl����2���s�B�if�'�W�$��*s⧂B�P<�$HfWT|�u��%�Exٔ�|���C֑_/���5G����:	5� ��L���9�䤎#���?rV!4� ��v��GP�F�Y�H����mC'xl��W_4��o����X���X���F�
/Y�}���
8��7_��W��G%��}h��D7�^�\B�'�\A��W|ۯe������,�y���"�њ썝ȇ���[,r}�Ӷ�D/e(��A�U���c�;W/�[m�<�G9��(���6�t�OR�h����߆
�7ذM0IxΩ�Q줸]�z���X�.����(�c�Aw�iD��'�������V�%��s,��r��U�*&�3u���iZ���p��֋Mw/,��j�}��e�e%��C5=�c+N*;��&L�WU��]~�Y�R�ι���۞�귋Q�)C'��L��!j�N<��������nG��A���n/�����"ڢ�F-��ٻ���.U�k�;�4�'��p����ю9�N>�A�{���R)��v����TI�?�2$�i�)~��7�=4 �9�w���#I�-o�����j�ޙ1��hE[�xaUTm��i����T�Z.��.�*[�!�.�O��Дs��Sk;����{�
�?j;^܆�nj�=�&�ǉI������695����� z"&٨��
��0u��dB�t]I�khw8����G��Q�wMK\�l8&؂ �5V�47�3��.3#Bp&E�Y�Gӧm��v~��
A�	��D��� �!ߞ�W[�����B�,��4���'��v��o͊��5�i��4�
�PgS���vU/ �1��p�lf6Ux�W5�U�b�k��F`?����&rrȈ��-4f�u�&�	��V:��D�h�dKΊ?�V_|ڋ�;ŻA��C{)����^y
��=5w����M�o����b@����^��vt��(��qK:#���͉ 9�y���:�g�0h���$6�K�9�'�v[���r����Wr܃��Y(�-�IA��c���ah/��X~����K��k<�n�i,��ښuT�����IU~j']�e�����񎾓>�HV�]TG-yU�ߘI��;��+ٚ�i��v�5�[�=�t�"�DB/49痔j=Y�9H%I�]%l/��DN��t)8u��u
P�w�����*I&�#!)Qp<�$�vi����G����]����0Ѳ#�g&z[��\ȍ"�Y����+��X��d�1���A�s���o����ãrnޓ�R�%334�L6e!k�a��F�r�P� +��Oc��w��sn�W�J/f�"Њ���<a����.g7���*�=�=���6%#R]� wG;����O�[��8ҏq��}cP	�?;���(e16ψ�v�T/�<"j�vq����6=�ڤ�	W� 8�����w'��wdPׁ������M�{7_k���u<���>�ʲ&/I�s�aa=�
]��V���r�)`�a�/UR��z/Ȱ@�>	?`�0G#�Q�.�#��۾ul%��Z�^Y�e�0�[�(�Ro#���י?6#/�#����v���$���e��X?C�*ٌ�@#K���U��&��,g8��I�u_��LL��,~
ƏI}l��g3����K�g2��P�[�hj[y��x��x�K]_e��������T�x`�����k|b�!�~��D�2�tb��Nq<v��f��wq�����1��o-,��w�����^���t���I�@av����Z�e	^����vM�C;��A�-������}̤����$CP���ϩ~N�5���$E�9(�>�qе3��,js�9	?�Q��^�� ��'��nO'Ӏ��Z��m89�Sv���W���2�l-C��Oj�!W���^�י�|h���+��+��tpN��k�IG��F?�Y�d�����QV\�JJ2�Vl�5��)>�w�������##�������Ș�	����?�;�-����|ը�ZS6����'Э�ܱ�[�r�{�{<�-0D��i��i�oS �M�� 
�t���������o�A&�*��vĽ{}V�����M �S��:�$?�e�R �)��]8Ѩ��1�k�m���*/XA�H�b[�\��x~�Ap-�]�Qv�.��_�9�(�h�NV%0$�,�m@����R~�ըMY`�V@ƪں\��@�
�ƪ����s~):h1��w�-��W���r��זzuߠ��gJH�	9j�+��)�N1 3f2f�m�w���.�&�
q\-��.��S,�qaq�g
@B�ʾp*�|���kpj�Ҽ����8M���e��G���w{��;[Ok�;(��V��$���(*O�3�M��#q�_��P�C�p��7�MR��&2&�W�Pn���隈��o���'/�t	�|�hJw�yZ��4Sf���F�pQY��c��*$妰K��6_�9u�����"���L7�*�/i�M2����y�ĘTL��ܠkP8Zc��d��
c��C�DI���l���6H�ˡ/�jVSKb���x�R&iձsy�j\��B�����{�}X������K�@R���C��g����;�}G�fc�CU�/[W���I3�C�:'D��_D���B��������Bi�N�i��I�V)�{�G��D�v�(����RoSp����Τqp�rp�;>�SL!��3��)��b1��ͷ���bw%I{t+����;p��������'�������fb�6�{p�:r�0�ĺ��3I�k�{a �Dm�� ��6k��_"և
^a�u'
�l�(���3`s�P����_�U?yf9�]X>�e%�#c��Ú�2�'���"ۨ��j��i��;�;͞&�s�R��k:��v�[�9��h��kgI��VBNd!��Nw�Ω�	���Z���yr�BL�ȹ�4(ǵ�ݼx���__6ɿ����;�C�o���U��O}�4[�%�l�Ae�z���IžT��'t�>g'磷v��}MczL<��c�`��u!��a���=M���cQ�m]% ò�f˅EHe���?d��hX����Wڂ����y5]� Hd�,j�����\��j���՞�g���p.��Š�=��]�?����?:��^&4H���w�d�Q�5�D��E�l��7 ��`���@��x�<'{.����A�޾b̬C���q�N�G�_�X�a�݀0���]�G�V}���骦���J7�t�yul$JU���/������a�I�D�-�پ�,��R4�m%�Ɠ�d�
��K����Z�A/��J}����8���=�����H�~��p�C��}���q�n"���g��M����]���aҐBt^�k ��P�����P�޷4��sR�����%��y��B����"�=,��q���f֚5(L���\�FM�*��Y􃶫Hl|n�}�;�Ee�.���w����{LU�� *��E�CS� ����B����өH�5" �͉�]|����@�n"r=S�D��'9f��Ѯ���N��E ����,l8���5,T�0L�Ӻ������ǈ
�$j��VZv�)� bv����������Z�w������kc�;�oYK�o�l�Ԣ����#]�����{,���(ΌcMs,y��$��B;��+Kj�9=1k ��{�­��ݥݫ΀�+ۊ�����tO	����i�#;K��!�k��4�d�Rg�+���K���z;�*��9:���r��@������d)��;C�W���M�s�9b́�FL���t+@'@�Bɬ�)748X��-C��`�H)����x�麀a;;��ӂE��/l�J�Z�F
J���^�^2T\��O�op��7�s�LR�s����? �7��-�e����h�Z��ᩔ;��q>ϘxVZZ|\�}}M�a�j��r���FT��۷� +�g�_��^Eõ�ݡ���<c��?�=��q��R����NOȅo�ř��?������?��K�p�#n�C��WpAяO��Xw��>t?�ņ���1�	�ť�K+{A�En^غ}Q?�޽�E�=�R5t�P�oG��7���?a�l�+ќ�� ,9:�=���w��L"D���h+��h8!�s�t&�;Zc�7�^�����C�GMp�D���z=�2D�9�J�tw�(m~���57�5���㌭�^�wC��˗*nx�}J8)-E`B!�Y(^�ƙ�l��l��Eҭ�V��n�x?�q�"�'ZJ��1��FLk�fD�<C�@�D�����?�4��h�LT^�5�BD��fq�s������@+�c�����b� "j�[aB�=���?��p�d��T��@ڢ�[ozғߊQ�o9zk:�nl��H���їZ�����-c$�ҿ�N�����'A#������4l
A㾎(@�1�ԈA�P1�2A�_���>��(�|u�'m����4Hb�n���L�����k�g�&d��O�j���z���'i������=8��#.u���1�z#�	��c�ȣ�5�SӞ�H��k �h�S��G�p�Y,�U賹 L��=]~��պ�5����"���ޛ߁ic���lLy�ƱXT5ҞF�BT ���5%��ۄ�8
VxAO5�f��[�����~���"������&�����y��1~�	,���@Z�!-Qf_g@�|F �7�l��y�qt{�<g3H���_�R:��65��+���T��[�Z��]�I<��+�D��㢗�6ب6� ���Nt�,xOS �.������b
/I��S��l�M���&��r�#�/���9�Xߋ�e|+P@>�;�Dc+Ep��1J5$�m� ���H_���OK�Z,�/p��B�\h ��Vh���LpXϫ!p���Rpw�
1�e����5k�dp^�3�gn[��n3uB�M��O����<%�1d���G���;��K#D�;R�~�~�/�34U �׊q�iX!L�A� H()�L+�_
/���~��cď�
�ӓ �O��e5�Q���ɻ{��c�����A�E�_�>����U'(���oQ�:3,�1�o��|t6窻�`�y��_���Z�6ʂe��}�n˘�>�5Ď|!����ai�hs���W��O���g� �-�c�����S�㶑'���
(��`��M(����%I֍t�|���C��3��Yw��~������5�l���S�'���|+��{'���nc��$����ce�G'�S����5�����G'o���v�����/Z��� �|��7�v���~3�B���c|f|�Q(1qB�q':��P�5�>G_��[�67Y������x�`7鳹FX��5']���m�Iʁy�Y��t��HW��*��!��?F�������dn`��c�T܀� P��0�����4b�M	O��H����+�ֿT�>i�Ox���ocl��>���o9諟�o�P�Q���2��V�6�������4ʷ��gh�|���&%f��{3�k�qd�oP��6H^��r7s��*ʅJ��}��{�s��y�.���?Q�#.����/���*_l�Ecjh���#B����@y\y���{���ci�ǋC��PU0Ah�ԯQ
��'a)8؋;�;o "��ؐlͦO.� �
è�mi� 竫Љ7)�^R�S�$�P�J��3�2�Ej�?v�q�����P��N.f'��n）��x`�������	���~hj-�|G]�c�/�˰|��.�Ogk �uь����US���~m:��hY�ђ_��z�j��a�l���X5�Z!��yw(��V������U��NS�>0&� ���ٗ=
��QR��!�>��-)6��MVU �j��jdf�� +�U����Yȳ<r��1S���{�-���\5 "�,B�g�HA��N�P�0b�x!��.;}�`A� c��hqy�t�Ե�@&�s���Ė���y(@�*4����|v�����>�6����0�
��������ar
iw�.{��G1��l8w�O�yd+���F�P ޑ�Mr�'��:��Q ޝ��h,���  s�q՞{?�9R"o�.mI?�+�T�����9����S���8F͟�S��G�\��F~P��)^��DD_�
��0\��������Y�Z�n\�R(N*։�Ϧ���gO�N8б02	�3tt1,�E��09��>! |�����W���&c��Y0��A&�#����#�������������{)�%k�=[L
�c::��B�or�1U�7�#i�ב����*P�		N�n��d�Ld�@ܾ֢���+���>b5��Q��ؤ�.P�<�����/��jhe8���ѫ�?�&d����I��}ۯ���������YЫ�me�e�.�`����-k���ʨ�it[_��+��l4��c�xi�O&�$���!�G�ǐA�W]��k�Cq���Fm�\��PRK� ��@uȟI�/�����2ЋRL��g�uL�6�H5�ʵ$�+��B�0���g0�k���l��?��U����1�1T�Ւ��7���\����9ɠ&�v�,#|Ye�u�,9����$��9)��"����6+tX��~ΞLI])Lf��S�`�xw��67�D��8�'�����MZ��/��)������V�S;E
����_k�	� �o&����x�v<\%~�uP����)�v'� ���85 ؕY�� PU����Gǖ)v��Q��1�&'��V�Ś'qi|��c���"��_~BE�0��.��t?����|��k�M8�@�Q~�M�9�ec�B��ꏩo1�t/C(nQ��tYb<"�fMד��z�>Wa�|�0�����/�6�ܙ��q�X�S��B1ǩg8N�(���;+��@�͎�W�����|pAǦ�$��i�-��0=tb1����d4ڏdL�B�#�����2�����]��R�3LPʗ�8���6�}����[\�T����e#�<�f�|�>'����'V�Ɋa-kO��2�������������eS�;��٨�1&N�#��3�����O�j��-Z퀬<�ڶ,#~��i���iJ?��8�1B�gvB���WIjM�79EU�X"���ɔ��ɮ�B��v��\�
��E�����nv�x� �TVey�W� 	�w�dƁ���
�^,���1����p05�Jپ58=�O�nHJ(��{����j�7���|����f4��Z�y�Lʃc�h�T��#�V,�+�!3�qsÕ�@>�M0�����~ћ�D�M��o5�s<8k [}9���م��~��I�>��ŉ�9����h�b/�@(���ʫ�8�`����r�;a�L��}Y !J�Q4	ԙwd�c�[0L�A�F�j���H��ey��l���y	���扉�U N�m��g V���9W?�oNτG)1`�zr�[Y5q3Kw��1�P�8���U�;iz7���-��4p��n�D��OQ��ϓ�:��L��Yple^;�Jhb� H����,�K��n-�j�� ��g�@^Y$��ZǞb�_���W<�b��2� h}��r��q���e<��AU7�}�T��m�ݵ�^�)2ղ��RM6�I4���W}��cu�s�wv�F=�F9r&9�OG�Rr�J��j`���6@0��)$2����5@>~�Y�V®��g\d�O�Z�A�I�B�uT�A}p*�\Գ~,��m��������Eh^�zÿ[U@Ywq��'r�@P	
�U@�m��O-��KH)d��"��$3)6Wn�2��v��}!��E�V$�@Y����hKrL�܄��a��گ�Rf�M�I�TxK��kY��n �*���b���0<�G�� �*��ͥ�}���N�7W�J4�sh����
ǃ�A��`䯅>e��*����L������r@x��X
�D�d%����[�2XL�7hpB�m�ɰ0|�
���aIw �C2�&vVtc��l���pI��$��NN��~¬E�	���e$�h�qt#h�^���[� vM���e�ź�+�)(��j�������Ʃ���5���i$0�3#�@�wQ�`�Y{�ϯ_��N�\����%�v�-�d_�����R�&�Gj��Oo����,�7���r>1H�t�Y���g{��M�dF��N��Ԛ!ǡ�<Sx�j]�d^yK�ڧ�!�u>�� ��4|�zN����u��V�%�	��y,@��kp�r��=��Fe�H91������|�Ϲp���5Dԁ��=�&{Y�g����<9"��(
m 8,t�H&��Lދv�]��p�jl�x�\v��|2=YW�6��z��" D��:D��O��R�F���}�����&\��2T�a�8�r�҂�2X���r�.*,��}�6���4�Y]@������Z�xqw��j��G��)�-�n50���|g9�B��^7p��4ӏXk_F��MG�tU=��ߨ�S�FƠk`�.�&�߻�Q$�����YQ"�r}4:��Q`����X�DZkx�jc	 ��ό]���fɑ4�iRD���8����UZ��6�i[��w��0g��"4ݲ�D#�J-O�%�'��lϯ�̞�pUEp�ďb�-��YT�B�{
��n�㙛]d����e!p�����d�*Hn��S��?�b���G�ƛ��
�(��H��.U�����R�*>�9�I�jޅSD�WB|s.47dW����T��fUvrt��JFҙg8�g�c=����Q�Q��+B�Ŏb���tJF�}�-����ܻZӪE���o>ۛ��I1�
QU������S���6BWB@j�����`S�o�����L��Q��lx"��h2�Q�z� k�@���)OYf�o�T���M�*��jTB�B;���Do���IH�Y(�NK	�yl0�ƻ�f��w�mG�0�L?r�Գ���#�òБ���$h�E6�:f�q����4n^�ᚇ"i���i�X�Y�M����sX��fҽO�[��-D�߭���\�޴ԍN�jkʅ?��w&,+��<�fJ�U�Y�>'�7W�w+	M�Eﹺ��8kV�?"�6��շ��N�Yŧ�2�*�{��i\td���_�=Ox�&�|�A��NYZF�����`v�~�R)�-EA�Ɲ���P*�y�t�꽠^�<x7�ٌ]�{{|�)i��`���'s���+�[��ko/�y�U�7ܰ�s0�}��y�Q�����}�	��ȥ�p;��#�ר����dj��x��w���&����PxƤ���N�U�����j*e-��*�;h������p�he��i� `�����}��Ү����+�X����,�K~P�R��N��Jt�˪�[Aop�Sh��r�j� x��|l�Qߕ�+)f�S�]��-���A�߬h�je�Jfr�/��UK��$|�1��n�'��o�$7.�H�@@Ĉ�*�V�=y=���GK�w�������	��92&?��ͤ���Cp�#ٵ�Ρbk�j�:���@C܈}0�U�<큦�*G�������ҵF���\;y�D��l�>����r~�+U��lmh�B�y=/0v��S�~f)�u�ԍF�0DRY:��,#]UJ�x�?��k[�������7��xG�em9q1M�_Q!4xb�hG!`:��1�E�s	u�O ����69<������n�6�=^L���,�}7A��2! �G.��+�Ӿ�w��'L��<ü�c?�3��ՙ���&+�ˬ��&_�Ũ"#%�lXs�ۙ>X��dqhK���5�U�/i3$h���O�N�b�*�Gpl�;��z:�S�_��F-M+:�qE$����Uxu��}�8��7nwGh�������.����}��0��TE��%�	����}X����9e��Q��m���v<��3y��/<���y�?��#�gGӜ�lby�p`��z!��]h�C�_��"G����ȏ��4U=��ɰ�7E�)%����2����-;���4/�g�r�Ɇ5��va���5��
)�y��+!D/b�oMC��������@�OKI���<c����(��l�p<)�l�,�3Q�a^�=��{�f���!'fkK��n��,��X}6LӑgI:��.�@U��S��OdMHu����D�Q�Ǫ]^<^c�;jۣ�P&C��	5�k�m�u�I���a�ö��6o�|�����] m�	���:NP���7B�Uo�z�U��s}I��ۀr��O��4<4�}S{�'�]�Dw(m�g��Yl��i���$�S�87�R2�;-���H/�Zڼ%�J�e'��衒�^���͗n�|[B,t��]�
�=�?:s��>��ٕX����~ۢ�Za�՘�1H�=��J>Q�\��������S�;4W^�<�&�m������x	�C%�x*����"���d��K)׵P�<����[�3'qW��<M����RA٧������9�f|"��x}2[�1Uc�4�@O3���,7:ͮ�cӨj�f��@9�u,u�#/{�J��rtYEpA؍�y�v#�%`�i	���Nɪ�WΓ��뗝�味[��W�|���L뷖�p=C�V6f��7Ҵt�N*�s� ً���V,�;I����J��1v�2���W��`�H9IAvj1���(�w�����^�����o�1�.x��kʛ�>���t�~>��E�������΂|����n�*R��Zb0O5����K�g�z��ܤ\�ۃ�b���,��n��yw����PT}���T !���:�cc�x,OD?�H�茬��E��g����@vQ��K�2ń���{Fr���mo�YvN���xQ���E���^��� ����3��#�gsA����	X���ok������-���>zy0l�#l[l���|�CEa|�Qr��X���~��F��	�?H���x���=��z�i�$��ӎ��9�e��f�(W_�������@��G���B�\i5=���cf�tBNA�jl�:�~�cl� 1�a�o���E6��/��W�������n��{2�&>��sv�`��~t�&[*��8!2"���-�6����Vk����8�6��$���2��Fi�k�i�s|G�p�Z�	��jq��d%��}b\���iLv�pRƸ�}(]��ϻ �U��i�<I5�h��/�@ʩ�����fx�k���@�δ�F���w����x$��������(ԯ��o?t����V���[}����z����,��D�+Pkf�Ρ���f����C���%�|Hl%��	����N�m���SQ�!����(2b�<�}v����;XP6��aUs/|����7)�hw*ոDi��~G����������2@Z���B�^�m?C�a�N�G�Ntw�����Fa�����̔��Y��X�P�����g=w#u��sG���D�Moi��^�G��g/]�W6E��:h�RG��!{k-k�s�r����h�P�����Bl�*���I�q�M���M��v�â@��ǐ��@���z��F�`��!^,�u:b��ݨ�,鰕N���l��H� :u��G��	_KTZ��{�v��6�������Y���U�~�[�x�O߇��,,��J-���t7����QVtb�����K�6"?c��)j������=���F�Ϲ��ّ5�Ra���q����r?���Z:5��7�&?0��x��������|�	�:}���r��+�IQ��0.Ҟ�E�fdb`Ϟ�*k�Ў���$��89��^(�@�wծ�"+`��5-3�7��ɣ�e 7��,���Q;A�2^��b1��ۯMq��׌a��7��{��4�
otB_
�J�ğ7�3!Cvg�˃kʐ��4#�H#��%���=?�|�+����n��ҹ}����djڱ�5�}b��Yi�wlD̒�A���n��.c�iQ�}K�.n�"��ʳi������nX2����-v��f�'������Y�>k�RL�O����O��<��k�l$Gx�p�$�%I����Q�hWe�/�?��P!�9�:O6����ڟOc�O3_�W�.$JS����*��}��뤶gs�8�w���L��2�n�9oRvŠ���:�3*�Mykә��:m?���2����:��Kĉ�o�}���իz-�t����L�W!�Њ�`�"\��_?k?!v "J�����9���1qN��k<��]�ZYA�r�v҅�*�}��Ft2ts1���8X����[��F����w��D��E4�uG�,�~�I&�����ƺ� ��Q���-oO���Ԅ�
����&�r�@�2�ȶ�{ri���k��E��p���u�s����t�+QS�s�X�
tޒ����R��b���h<f��5�^�{+��RX-j�Z�su-�J�K0¦0���m>�yQ��?i;��!�����4�J��u[_��s�C�~_G�yM��
�%)��N���c̈`Yf�w�������֝��[�q�S�!1g�}�Ҽ�z��3��?;�B����iT�1-�$����D�y�f��F�F�����������Gw�W�H���i�x���Wj�9N���������S󐀭M�V��I�����ݢ�i�aQ�d12�]�M��K�D�@����^��`��csq�� -�6 �e��:-�z����� s�Z��-�X�Y=b�E-���5�++��?����Z+�)��	Wh >�y&��O�&�����J��t��T����>J��#�*� ��v��s�C�[Ֆ&t�o�;�%��vߕ�}�Č#<�(��8f��V-A��h3��_]>�wm��S1�:�+� �\��
�;�:��&fSq�b͗w�_/a���pBŌN���J���'h��˸�C�(�,�ƌܤ O�p ̽w�EO�J��K��0�}Ď/{z�%=T����}�t0Q��K�_Ͷ�� ��̤��#�k�!#o|���Q�In7v��/Ƭw�?�80�1oR�jR�q�h��,�u�}˸��7�������"s�z��� EUXOv�Q�K#�Ӟ�n� �&Q�����i�з)�yEҗ��sb��	��Fǈ!���N
���ya���6���P�8��{�Ǖ�Jx�o��3�(����[U	�`f�q��⠇��h���DpT �?m"~�9*ު/�-�ؗ�A��5��uI��%j�ݜbI|H���������6��6]`vw_e'm~���ۯ�~����l����yj�Z���aN���9}u��K({���{5C[_|�@��V�˨6�����H���:����l��P��D�z�L�?JǠ��r:�h��?�n�l�Ѝ�}'� ��F��8q� P�e�W/��%��I�'�]
�6��6�A��Ԡ-}���=�g������dԙ>KSP�G~5�s���OY��!��t8P�~m��ŧ�q#�lЀ��jڟ5oF�Ο����qq���z�u)a���To��y��)eo��N�xn���R��箖��mᆷ��x���Ta��=)׋�I���c�ӄ��O��DD��\CZn�XXi����6%�߲ap-m gZK)���5(�!�s���b_���Ъ�w�f���U$�3C/����k���(�հ{:	�7EZ���� ��<�_�S��9��&����<�!��}� ���}�X3D����d�K=Hy_C���c�_O���$3d����o�#�$5��Y5�	������5�O��`�&PS)���V�;#��ݧ���5u�K��~�=�7!�?I�m|y:�q�߭���_�����V������(�a��w�e���p��z[J�a�7Ǜ�5s�=�9�n�(�"W��J�h�?�;0�$x0Lu�R�Y��
T��� UE�i)�}��'������^:�L2�X �+�e�2�`ؘ��=u�/�i��N�ԂG��Hݬ��W������~{��҈��(*�׾���������1��T�������s��T��ޓp���2���^�?�h&hզG�7�2?y*���G��5����g�����8~��UĨ��"� 	9)���\�%��`7v��-N����(�f�؁���~S����q)����|�r{߇U��U�@:DPR�j��=H�P2C�J�H�����PC����C����<��?[��?��r��u�u�+���Z��I��x^a5d�R.R��%��m99[�.���a���a;�6p���	UUE��)�.<��`4��OS)@5�4��P�_o̩�ʥ4 �^����<���v�rX1�����53���zC��n����{sxn&��@�s
v��;Z^���j��ɺ2�K�����7�����E���F-����j$��u��	�6AY��t):����t�������RJN}��pq��?]7����|�vc>g�ťiN�O��_���Ͱ�a����RǓD���q39����y�pŔ����Q��j��d��H��K�ȏ�DSL�c���]�����C1������}?��-=^����wQ�q��ﬠ�G����2F�!*C��ZB�X$�Gײ�Mm�YfWr <k ��~亷d��any)@�U��evR��o���	�}�,,'9��R������tuK�R�w!�/�/(-����,34F���B.fW�$C�?�T�M8� 1.�
�I8{7�;��CI/ז���7-�u�ɗn��Km}�?h� BI�|��hcV5�Kqa��V=��?x2pR�Dr���=��0�иjL����Y������ň�T; ��6�ƿ��
\P��3
�++�cu}��x�7bQ1[@�-lU`��o��'�:����+��v-��	;���'m�Z��~S���16ߺW�*;,<�k�˱�$������~?s��M�Gw���R����rt�.�Ykv좪�9���t :�������4��^�&
�bt���|���b8����kH���K��Q�9��<�;�i�<t�#.���L�pT'��x�Ԯj�9J������!��#@=WjqsR�36ˡ�[��QߣU���4C�OK���ҷ�_0����DØ
bX�0�͗���S�}9��6m8%}rm��(�<���dm�WX���Ƒ1A�Z^�4��}�̤�� &���UI��E�D~����n�;ڴ���)�0��m3�`�ۜ��D��R�(��uuX�^�4Ɲ�����Z~��I�m��z[e��ӽCt*N��-S]�Ṣw�ؕ=B��f�����*�c���e��7bv�\���>�ڌ�2��
za:���o^�����;U1�8o�bnCJ��j�0���������3��W��*D(z�c��h����n�d+"���1�y���M�'��]��ge�9�9�8���>3�q���B��6o^�y��^in)�����r�>M�bb�� D�KNK��;j�6��������^�h��Tl3ˋ��9��� x��`��f����*5pQi5��ќ�������>��S}nG[���$�:���k z? �?�L�tP%\��jY=���],�t�c~ߢ��sQħM}C�Uj��U��@c9(�4�5�9��ҳ�t���`�^ˌ^r��ǟ%��_|�6��+��{/���p栱��̐���SCaA�F܌��>�Y�L��?.��ќY?��Y4iq�b-�'m�򭬱���^���s��n����Z�r�\V�XF9�<jh�C� *ol���]�WR�u��(Jw77���G����~0ǓLe��v��(s,����-��ƘYi�D�ѡ�B��jox��? ���y����4d��{��(��i��Ծ��$�r��1�'�?}���p�JF,�����r�d8���[$�~W�̑gI�3�|{�̗0��~�������G����{����F{U*#��0U�)��up�*M�@�Z�F��!3>�0-+��:j�0����ƙc�z������+�n���ueRq�}�
=yt� ��j���7#�B��I��(�J�;
'�٣I��N	E��:3U�x���<>ʼ�#�S��C�c�R2�Kp}��Z��b��E㴇@.�S�S�q�����M(L�e��F`��Z��8Z�㗥d@��F��M�	g�CXsl>�_���j>������is��'�(��Z����H����̙��ɪ@ã��&�-�n��H���b!�]91g�[�}����$�Y�xA����Wv(.;�:��J?n	:���ز��BEF�� ~����I%���`�m�6��w"�d�6��8�d��o�NohY����oTXgϞ��:P>�P%X������ՙ�-3!�A��3vv!}���BTqXpv�kkcc�U"����5�5����Óڍ��r���=��5�=\K����Q��ꁊ���ml^�ЯS�>��L�E��&J������Z$�mW�,�����5�������FTg�2��rg��㩽��ӮH� ��*6(.���)�u�p~���R|X�{P��KC�h�B�ڌ?Yd]N��5�Rs���1�:t�����2z��t����0.���eaJk������h���k�CP~�P���;���_im�%��&`��?�J*�_$m�+������J�k��������Ҹ��w��}�������ؐ�D��ٳy�Cq�@Ъ}A�3�C�+m��ƅҬ�HPX[�"~�F�m���e�Jf&�\��PGyee6���r��ܲ���Q��%�*�O�ٟ'�t����a}jo��L�^��nS���5�Y�-�㼭~Hv�O���[ǅ��H�o��L���jr�ϖ�n|<Iw����}�6y@p;�:;�˟��d	�>�I��V��������9bA�Ж�]�㤫l���\@˨��m�C�.��Z�����|p��eiOܤ���� 
���w�q� �y��I,���J�ge���s��@v��ٛQ����-�oE΍�J�̻�~������f����AB�3��6v�V�#
��їt�1�i�Bx7{��s�{��j��A P�	5�	��{��ך�����7��\�'�����囗;���X��"�Wm�~E_#��>I���<P��xM������@R��oM��'%ȋ�į�� M��/}IQ�m%{�ѯ"����`��t����2����d���i�q_�Β@�p�V��݃����.��b̷qtmz�> YOEb�
Z�!ӭ���J[����C����@o�I�����d�9_�l����I��G������7�82
�#�f������S��ɀ��9 3@�h��o�r03?{�|���'
��r #{�>�$ܱ�A��tT�W��U�	3'�C!VB�d�>�����w�ߚ��F.�7R�[`��l�|m�?����<{m��<�o�
���N	�Γ���~�q6���eitߦ�ƏcF=�p���7?����n�O�a���|�g��`Yj�բ1���7ۏ<����;WP�+K�������v�Z�#�UBr	(ҟ����xӍf��틓E.N��aޥD�s�1�t@��������i4i�'&�?��ڿ�vT���9Zn5pp��^&�)-�h�����[�v/X���W2�??�Os=2?��d�m��c�,s��Jp����rxYFs�CKk�,��^�..v�sΟ���S"eP�V�c�a�^ �A� ը�'�fɉ#;J��{�_�\9��-VZF>��Nc��H���&�ƳQy!�i�BB���qc��J՚u���XZ�l]�m_�wH�|�jG
��I�g���	I8��:�8����e������#x��Z�8Y�z�Q�8����l)�a��]Dq�{�x��~Lub38�U����~EV���!�8*��R4i�hk���֛_��}��9�8�b/�� X3�%�sDO��������.�j�&��]����u�ܣ��O����a�~$F�`RKdl�����sn':�"uZ�|'�̩�;��}��5�j�-��f7�
^i�������hXc���h�h&���J���t��-d�u�'�R{m#D���r8�s����%��2vG�%;B�t���r+�ۨju;�
فW���u`jF�N&��gC��T
��>�`��;��SOl�j�k�6������0����0J������H�+b�Ϡo_��c��9�U��Uo��L�Ԯ�U<S7>�o�O]K������Uà�
�Z�StN�m~;$�N���>2w5��`��2�S�;��V��kO��������&Ǻ;So�����w�Jɹ#��i5�a��}���,JQ�2����H*n�#v�),Y�&��+�>�������	v�Ǐ[�mY�"�I9|�WD���B#s��]+���>j��#��f}R8@T�W?�,,H%�#z��N���_~/�]��z���.��\��D�G�a:�g�tp\��	UU��%2�O�+�]�LJ'��t����M+�W��tU��Z�� ���4��'��
.9,�fcXS)������Υ�G�+��hKQڞ�GU���������_鹧ߏb���4A�t��5J=+��T�hO�ɼ�_�)�����U�;#�ú��E��'�A����q3=����{�0#L}�a�Ѻ�X�Pp��$]�j�y@{���ll��M(�&s�]Q��޼"_4�=�1Ax�`�im��6<�+Hnv���,�G��2�[?���~���Jo� �i�twU�F�]�_I�A�KջY8��W��NU�5M�<���Z���|f��43�7���<�b�~F����&�-LѪ~N��>8�s���X����K_JxIߨ͸��'�&g���퐑#;vy�����.�J�Ne��#glW�{yWww��b��v���`�{В�����eS�m)h�v���r�{�b�΋r˩�d�a��������N��zf�rW<N�{����k)�J���������n�^�t ����ś;�E���+S�N}�c}������WL�ο�y���:EqmH�=�	�(���iv��A��ۉ������\ҎC�(�ra�N�� ����;����?/�9�qb���pW�Q��ж��3=9��6�\����^̳��(���ƣ���|�;���
���=J]�W;��~B��_�����S������u��Q���f�y}��hy~u��m�vQ�ڱ�=<L��C���Z��	���䉄�h�p+�k�O@�t��|�J%�0�jC�h-f�����B3������'�1y�e��/:JXfe��Iڥ�b�i�;�l��&jT��D|�S����ou�z�/����3V�n��@`�Wwk���:"�j�3M��5�^�j��ٙ��ێ�A/�#�l�ޑD`��*aJ;���7q�9�T�n�a�ݙ������6��)��d���2��v�d��iG��S�;�H4�ov~T�KV�禝�G�����;Ny4r��:��eW�!\?,\�VQ��<q�
L.3im��[�����G9ĥ��\���Ҡ�ɡ%	�I�%�Rt�@���$4Q���ᰮ�������h�0���xs��p"14/ ��(8}2���/�R�����C� ��t�S��X==�(��ld����ʺ�6�Z�A�s�_J��I]�Jz�(K����;�����
�S��'Q9��0ԓ2E{�z����/��㦜<��	Ykw<C��f�ײ��%A�q;�J.�g1�I��>��rQ肸�r� 4��,;j�ś=f�3꣊��1���tϦ#S�.ˍ�P��DC���e��<a°��d~����1�Ҽ��]	+b��Yut�U�cB�V�O�v�/n�{e��<{[P��������N}t��U���b��/%c��x�A�ÐddL}��pF�L[#6&�e8��5��a�9�5��T;�/X���.>rs�j��Z���Sk%�%���p�Þ�{�s��#�u�Jww��2��?�	�q�d�ƺϕ�������>���U�ب_,�m���6+�P-�v�'Hr������&h��5�%��ٺq�1:@�p_P��Z�D{l��� �VK�{~Z]�=�.hZ�U-�29����Zp;:�۶�]�>ԙ��8�`h�����Wj^96�9����#uB�E��,Ѭrf�FH�3r���5=�� 2֚�N��e�f�����(�i��pֵ�Z��{/P%���K�v�����W7YmY�6����c3s�<��׿�.:�+�>�u��l$�W�i�Mz�1U�E�є#���gd�Jj�^hUo���Ml�W�<�P�����C���Q�8��ķ��tbr,uU����D>ډg��2$p�Z���Ƣ�� ���sV)8:�����GN��E��:,���0ܺ3�L������C��W��@>���6zrX����*���t���Gk�U`���c�W��X�"�qku9y[&U�]���1�7���A%JY���F��=u����у�g�YV졣`�c��Ȅ}��t4�Z��r >��A��bz�D��
N�`�� ����F�cjq��J,��U�e���u��n���5������^*	�������8Qch�����8���y���~Ƚ�+��ߪ���<��2м�L(
�z�H�S���<&A\���^ܒ'"�e���rx����˯�q���S������0}�46��|��r	�mP8�gc�^㮘nT�DV�+ɕ/Jh:�N�I�9(��{�H������,n0�<�Qv�Sv���^�_�� ��=�ɉ�B��U*ģz�@a��`?����o�82��_���wX�g�I�E~Ɉ@v�A6
�+ lD�_�p�]Y�VY��"��jb^���tKk͝�\1��"t�3^�Ɯ}�����-�yA��}/k��U�
�jy���'zb�z��}Q���p��{�ޮ��a���yi��$�O�mY�%}�@�Bz�PQ��������
��Z�|��)|��t�����GAj�Y�䏰]�W�S�B���l9V~�O�&�w_��k ��Q	/�uc+L^�|m�ž-ܚ��@�����뤖�urs��;l�!w�b.�	��?C��e����1֩h���k�hG7ӂ7��^�g�Ld�=͗k�#l���8c�(��
C�m7�@v��&ʀ����ڻU��n 
$������kn�a�DOH��J��޳1��"�U��L��j�s���m����Y,��Ve|g �>,�bN�K�8�K�G?�x���q5���r��-+&��J�=�-�v)ﯨ��m����[�z҈�JأlP���,��j��X�"vKZ����6�t����V�����V�C^�X�}`�����Dll�ܤ�X��2Dv����02|!ۑ+B�Gv��r���\��v��u�v��S9�K��oS�)g޽|��o?S7�ܔ� �[�5�ؐ� 2�lm���#ųGz͊"�`����[@QZg���q��3�"��C�
(�K��/y{a+v����XGܞ ������s�6-��1�/�̴��#<��6�l��*}������`�?������~���q�Hz?��0�m�˸'��Y�I�'u����ܑ�{Q�X���n�<h�d��6������Q}	*����wgC��4NP��9s��S�n΄`�9 v�Oa'��������\:�������U7q���-O��^+� �^�U��1hg��)}��9��~��=6��'T�/��~�-�(�RX���m{?r��\e���콻e����ޙh�Lg����j����vkc�=���g�5֊�*`ĕΛ�)��8WL������r���_r>��n����)ޫ	1��w;?�����;ͳ���H�R��ކz�"Q��Ѿ��C�,d_sC�D�+0O}O��U:�<�]���u?�ȝzXEۦx��K�x3��������!?ii˨�<�	��=�F;�����2.���T�c�$�JoH|T�sT�*��=ڗlx�ͬ�H�u5[���S�kӬ��>�Ud������ّf�q a3T�U0�:�Qa��-AL0���O�	���u�<��98�UȎR�a/�ۇ���ȷJ,���3U:d���RyE �� V�%�Z���]�y�Y�w�JtP�6�̊�D8�=�>��L�s�$�Q߂*F&�v�1��k�0-�X�x�7r$���+g"��F��R��������7_��Lq9IO/�?��Uɾ�=X��ZȒX�oZ��l���U��1����&]Gs�&�4� �GOI�/oAHE�Z��U��E�.����a��UU��9 Bx�,oi���b�X���aB���K(����9�óR���Z�uX�q��,-�C�e���o�R�M�sT��W�W��al����`G1/�x�@��� �3��7�S�(0=��[So,N~p�Ʊ$���Uu�au���^�# �c��r#� ���g���z|b	3���j���J:(0�R	7�,Y����gu7��Cg@��CE�K=6%�����V�޸2���S�q\>r�	�;���l5�UspZ��Ϫ�ᴤ�?�i��B��h�m"����!�Қ����	���ڍ���H�o�3E�����k ��y%�_��P�@lV�@e��]/��#�pX��rQ}���	��0t.n��!H/�k�$�}��)�1G��sD���9�C'j��B ��g�C؆���[�	*^N��?��Mw`K�U)P��A)( 1y����0Snk�{{��#�"�7,�%��}Pŭ~�#hm�ޞt�f%h�,�/������c<>suIC}����%�����A�4��>�c���e�+C��<7��/��)���aH�{A#G�%)Z���?�q1�U��G�Ǡt�*��ꘕT����댏��lT� ���<'�a��K�*�U���� ����"[�P���`�٥+iA����g��zť���G��%9�e��T�N�e=@9�]01�?��N�)����9�$8����"��-k�����������)?5�}�li����D���7M@�������ω��\g�-��+���V��.aH����N�Ɉ'a����R�m�����Ge-b)�̔�jM-�ǹ~+�"_�ja��C �;=��-���a�g�l��^����S��*�dJ�=z�H�����X�b��^��+�N���F��'�p���=Ʃ�&�%�b���͹���-E��]<��5�ҙ��>I��ӯZu���M�^6~6�2i��%�p��B�$p����Se�|�	��4�������� �T�;�H�ة~����W���U
�z3�P��#���IB	�7��
5ֶ�Vmv�Toa���c�#��55ϖ;7��v� f�'��9!�Fb�G]�@�)��d�3;�֡���e�N$	5=��m�Wܝ3S����65��44y9Ǜ4m�9f�=b#W�&��[�DUo
c�7�+SP�h��k[���y�>�H�΄��K�Y-
���n[�?���e -�-�^I�Gҷ�i�ѦǣPq�u�}r��=��D����n�?�uKW�8ӻ�ɚ����� �֠���6���J"P���Ƌ�M�-Q���W��9crΧi� =�:��=���� �('�_��C7�� ���@'���E�ͱ n��h�{p�/�r=��ΏO�x��; �] �v��u�8U!��kՎ�l8a$1���L~A�C��q=6�~F�z����;��b��񦣮��Фw �Uֲ��q#o�Z�ڿ�  	�죊m�vP	7���)6S���sG�V�����T��=�WV� ������1D�;�h�>���Y@�%��S B�>/,�HE��!�{w}uGΠ�A1�L�%��P;���E�4vTB���g�-1��/ø���%�gQ���&c&�M�}6�5/���|tF�O���M@�p�T�0��#�=�&�(�W菔�r�KOL���23b�!l�%���k!����pkk�]�f�#�]������x�v��A<^?%�o#����D�j������U81g�>�Һ��ӧ�����Kz���Y ��zڲɭ�9�$'�u�ՌU/Ů�{�� BTug�A�cEI���x�"����Ȩ��p�����U���0�|��̱��N��y�����nІ��X`'����^`츷�P�I���v�������(�?��܌Ֆ���zl�>֫�t�1۴.l@���t����Ð�/��f�ӆ�u�����8׎W}�>z����|�n��7�osR�+w��u�}���k���n�BZ��qmp�*!�H[���еfb<�<������1��s�]�{i�K>��EG��G��;s�5Osy ��k)��q|�񹀢 ]�P���0��Y��G}ڐc?@������H��H����� ��|�z�m2m`�]w����
���Nl�Cm>����7��,���/.,��Q�it��3��Ν���b~���U��pk�5��D-3O�ak_O�-�gQ ��$,��a�/f M����� NV8���GPIwTMʡ��Z_U��.7���R�1 Y]�[e�Ic�1�04��5}����K�:��Le�gl%�}��[<�i����?\��? �R�Պ�j�{B���@g7�y֯������/�˫�)�;t�Bވ���l�zCG�[T �R��m��7�`X�%'���B虫��;�)�����>��K��f7v��Z��ǘp��y����������j������7�����e�%�^e�	ꣿ�}^UR��� ��ky�<�_	��i5e�H��ȗ9密���S2 ����qmq�˹lPx�L�顊 �._hlx7���Ўn]�2+v��[,�Kj۾�������>u��A Q�_|���NFp�V|�t�E����+�_®�� dC��8��� ����ƍ�u-<Ѩ�y��qyme�ǉй�?��no:	����8�!�u=��Е�&5{H,`��c������O���j��T�=<�H��Irlٓ	�#����I��FS�%�aP��5��4솩q�:��B�7���D�L�_X �xT�S�Wz�o���Hۜ�$��~�#�Cn�*�Y���`ϯѠSfs-�2.���"L��E������d!�C�v�fs�t�Y1�e�v���G��T��J�'�d����+�;P�ML�>�ո8��q�t)�ؙ�X'H����F�5ޣ��ӭ�� :�,y��u�@���x�@�!O�y�� �f�Ʀ⌕0�{�#[����6XA
q���yg�>o�CO����x�`������
�?�|�"�Qv���-n 6�9��_9�+�2��V͈� ,&%L<f,��Ɩ���#�&\;ʅ6��*��	ӟS�O,��1���V����L{Be�����7������E@lx�a%��>V#+�G�ih[�)���g����
���7�3V���ҟf���}�L�ͭ
s"���mM�D���@��K���s/�a�|�9�����I����J0޼e���w�r��p�?��h�u��Tfp_é��+��>4v��_��]�6�q,�6˲/��s��##G��ja�E�5_���_�,�%5���~����Ā� �Ta��\8�i#�n���&�a�@�}��^qN�8��K-!���+�����i��fwD�A�*O�4>a>x�f!s�Q���9P"B�`��޿e�-a����$�i:���=-J���ڡÐ�7_M���D�6&Ѕz��(L��7�Պ�@F�u�\M=���ގz��(GH��M�D����uϽx�ޤ�*r�)�ԇa�S�Mf~F�������+SyqQ��)Yh�5Өw�6�����bS;���R�b�8N!0���t}��+�:H�;���n�V�II�=%gwٍ�qߺ��xI"�F����s�O�E�Mp1mj�*��^�O��l���q[ Ȅ�Y-�pT�+/\C5R4��2YV��7��*Ӵ����ޜK�&$%k'�l��Y��{_��[}��\܌_�* ������7ƤL��`��@�{z:��@0�߷��R����b��Dך�՝�O�h~���,qmZ����譩�)�r�֦A�a��9(�@ͣ�Wl!��y��s< �#e[�N_fLP��Ֆ�Y-�wb�uE��i���O�kH"�z�S��|�<��@��f�)�w�a�-�A@�u�0��t�sC&�6�+���l6��g��%��쒌�,
��>(�!����SS!��q���YtSq2p?���z�_�G�+�^O}hП�|#eЙ��؃*�M>��JB��S>�}�_6n^�˨�|Gߝe<�7� ���Ạ[��'�r��C�f�J�i¬c� ��,z�ƐY%���X�3�?�ޤ@ߞ.�z$P1%�?��	��bH���E93�P_ a����v#����H|��1'�j���RJ'4Ԙ=W�r5�u�
6��.�K���K���Sl�y�c>���5���{�>�Uy�5�Z�x������܈�OjGz�0���G}����*i�Ɲ^t�� ��L�og���+~P��h�>{���m״{'�����L�œ;�V��������Oj���A����jW�D�[��\s����,|� �����iw��V�`D���z�Y��2Ґ�6�aa3��6��Fǅ\W���zTt-�t�`�\f��0�J����{DY�p�)��|�H��{2�,5���*�6��\�m���nCe慨�0������!�]��h�S�d*i����8�O��T�]�>,̨-l�͊O�z6�����++��;�N�V�-%q��'���|�:��b߿5�14��'݈+�t�I��#m�u'�Z6��vã�	���,�ukE�N�d&�����Mq�A;�*�i�|T�2r��ϝ�5�h�����m<?�T-�Ƀ��.�N1�"�S�C>���h��L�Xǲ����(��b$�z�s �U�y,�1�7>C���w�R���Љq�u'B/�,~��ɌC���`����YF�����<�
������m��Of��͙wY&�i,�.RW�0EC3!����_��sZR�
�j .� �z�L�{ڟ�1����_X��öh�\�L�a4���,#�*ؽ�>{K�G�Dy{�rj���Y	 `/�pA�������aP>u�ʞ���_�:���0��ֿ�&}Ҵ]#'mk�92��/��ND�isg��b��\'�$�y��w�-͉�M�u��	��r���Wi�5>�~l�}������ =�����=�?M�AB���.�hq(�n7Ɂ�l�Lnم����l�	��%$g&d�@>B�����̛�C�����#��ߗkM3��c�>f�	s�5�<o�Z�oi�����:Ǯ#������.C�Cέ2��@������u�+���*��f:uȕ�J�35#R�"3f���]�{� �o$��N;��Ƶsȃ.�+_̿aDB�X�%���Tx�݌C_���2����|[�X�����K5�NX��x�M���V�W%������{�_e}z	���JJ�o��P���S�XȔ� Lru*=��f�����E��\��<�.BPAOd6ĩ>ͫUGS9����m�윟�X�[(�"�Wf�F~K�p'1Į�����c�M$�����M���+&má-nB%���c�_BGx��m���xk�8����A�$���{���e����J�����lw�/8��w*Vn�{A��'��o�M���T"~R�:%u�Q�M�V�+SM:��<sR,s�w����p;�+2+e��3藏���@�-� '�9de]�C2���J^Ss��� PM<Tp�U-50};(���霒+wR4��G:� �lbd���Ξ�}p��������ʤ1�h�Z���EAR�>��n�=�C�����@0�� _ă�'�����Pԃ�M��_�6�
�olU�ݏlN�3"�$Q��YW�@�����&����2~Q4��!L��QO��(�c�ȧk&�c�r8-��c>3�%u��>�X6+�8����%��D[��W�E��pR�"Eb��2�)�@�MG�wˊ��6C�4�7C�� �����u�)X���(� �l��C�����dY���zR��r9(��(ě͊�v�w�Ǧ=�	E�'�yC/�� (��+(�-F|B����F�-����j$�|j��y
U�[0����T��PZ�H�P>z�q�t�T�:�m��q6'�bˑ�o/>jT�P��3mT�P�W��_YLS��m-�}�-1J:߁�}͝M��A�.�x���^d��z�ⓝ�f5�H��Wyo���.._˥
2Ɂgr��Hp�e���4���~�~"��7ϗ1���$���6�H@��SD��3��{�I�Y�R�^� Y����'�@W��"&vڅ}�u�`�P��l�%�=1A�#�_���+J���;7Q�]�ꉤnV������Y��E魊h�.�*��*�1���xmg�ك�w�a)n����u�Jr�+����k:TIOm�-"����x�qs���x��|�B��퀊�J���JA���a���r�>/h�b�ӕLd�HPQʅ�Y�^!E.��lc׎椴X��D�,dG(y��s�A	�PSU��o&A5�.c����|��T�MZ��� ���@�|�v̎�ޞ�5c�ʙ����?U��nc�$Lʒj,��(�z�N+'�t�+n����H,�<��A��#Z^�}�YG	O��]٤U,bpoN��D$�6�X��**ߑQk1��֚o�\\��p�n���+��.k�h�ݺ���Jmʷ�gֿ�Eɧ�����I�=�� @�C	�����q��<���87\���.��6�iP�=�	%��Uk��Z��^��=��*�c�H����1g��nZ��b�ܞ��T�֔%���3�h���<��	�44ΐ��J���wD=��/��U�~���FjqF���б恲��=�h��=��'��Dw���g�O�E�K�u��V�]�*�:��UUq!��~P���Ae���fH?V��.�R�o�k���nPO4e��F��3��Ҍ��²��/��iy���U�������8�;���-�#́ܵ�g�b�cE�ɦu�����A�
H�=@bS~�_Þ��P�w��;|kS��n|L�%TZ�M,s5]4��Dg�n_�d	cG�i{�Dﺭ�śv�K+1l-�H���&�86'�'���l�U�w�>(5W�2�:팷�19�h����#��A�S���~��NxR������+����D�x�V�K�%�NnǶ1��&��a�ea{b��!L�|�G��יp���V�v�ϵYo<z��~��e`��Y3��4V:��1�*�N��zـ��)[6Q�}�\dS�V�wK�~ӎ�x2�MWeA�c����M�x	1J���`��jqr�Γ���xL�xD$!4��{̧�Q�I䞆���|����F~$L��1h�z������帏�^��s����ٹ��޾��Cњ}�1/��*���Z��� #���5z�����5cw��ʴ;��4ua�5ջO�Ƅ���L%�I��bvT���$�v�]����^-���.�AfY����g�Y�4���=�7'%�L�E���ZDD�M6�R�*�2� 5���$Oa��a������ʫM�F���SDC}"����B�݁��ƞ�����s�<��~���8�7;;���W��_'�F/�З�F};C�L*��DB��_r������9���c1o�4-���
n'kk{�ˈ�փYN�Y�"��f�?B5os7�w�z�2��9��Y5 �4���B�<�� ��K���MZ�*)��<��D�|�<r�]$<hR��w�jړ�\��t�T"�ʛW�y˧�:��/��W@	��{��PLa�������F��6��1۔���J/+~/e%;�������j��1����A��0�Kƅۘ�k�W�&4Ǉ�ǳ�k�v��]b���@
R_��a�=Wfq`T�a3�����ڣ�* ��]O���������>����M�Z{�N8�"=e.��}"y�����U7��i�N����l�.�C�Y׽����j�����vQ��#/���:<���(P5Ӊ>�u�|��C�ﶪ����hi>�	�^�\�� ����Y�}��9�Z1f�_��-�h�a^�^q�%�,� ����٭���ۯQ�13�86W�E7�����@�#(�1�B�*�L�o��p�)�]��4���Xt\��������,�0�p8�C]>v'_��]������	�*9�ɛ'H��&������rݐ���Oi1�8ݗ]��#Z7��7Q�]��_����*�=Һ��.�2�^�=7w�@6˗K�s�ZF_�2x�֓P��c�Ly��ٷ1��{���S���a`����oh�+#������Xޒ<��)f�����[�`-�q���*�j*�1<C�jFNU` ��e�ݔ�C%J������̎Kz�������ߤ>o0FE=�Ѕ�M̓=��������k�S�@�ny
�F�(� Y.=/�{���o�i`�
�q�$�
+�%w���K��V�#@�Чګ���2o�F��{��M��c���'��O��*�=]$ʭ�wd�i�F6]����[�eWo�f��p�䤮�~!��O�|=��$k�U˗�^˝6��TP���w$F�v\����`z��B��Qߞ��Z���L�3]U�i@��ϗB|��N46�z��x7R�>��k_޶�r`������4�1�G����)���Iqu�N3����)Q�	���g�)�|�tSO��۷�_K&V�3�I�������U͡��XQC�
���~��S�z���q(��_�
�g�5����5��O|���R�!�ĕ��!���]���d`��ӫ�(����B˖�����qÄ�
��L�g3���y�~*��*��=a�K�9[�Yr���gu��K�=7EO<����V��6`|���PN�J�g�"�%��OA�N��1��Ҡ7���t���!��:d�+��->T�R�ĭn���L��~׭�jY���D�6w�}���!����$Wh�1���h���VJ�W�5A*򜫑�>��w(�=ne�rw;����-���)�rC���׾���ۊ�([��0}�F�ޛ� �֢���>,���i�f[���"������Q�-
DY�ɍ��� �w�YW��~������&�$�4��Ic}N���x�u��,�ՇF��Z���Tp'�m�1�<��{:�v���6��-�����ʢd6L�G2(��b'��xl������8ϟ�W��:[���g��pn���*�P(��=i�f�n�W<����iC���|���)�nf�o˦� ���zR�s�~bc�G�m����<���@�c'����PQ����(~U�ŠCI��i����!�r]���D��A���n$fFrh��g�����=z���{�{�s�[�w�B�SQ��ϯT�;�C #����	�u�`1L���w���T��u�n��s����JH���VM�
�P��HA��>��7L��\_�6u�A�k����]��R�E��p��P�����̕Ŀ~,ps�[j���̷be�~p��^�]w��sTׁ���{ޠ��D#ؖ�[�M��U[�D�þ�oe�~<�M��c��!F��p�e��'���lTǭ��8�����9-qr!Ի�ί�`T7�\`�sw6�>dT�g��}1){��f!-��!G�d����-��	�yFj���\�����d��Φ}�OU4�aS�5�VF�dl�"���F���͎ٗ
7 �~�B���~R�_�\�q�?����!�q��������R��NZ�����nv�v��u�6��||�F�;<�_�}��J���Kum�#s�P����o��Ώ������EҖ��m��F��5�0^�Z��;?�����C�4ee���^ca)a�-(����
�>��x:j�"���:�(�$�In+���2�������?����J<�5��~�_d�c���0��m�����c˹�2*U������U,AXZ�/3j�PݵIV�V������˿��z�B�=��?R�o��'�1���x��V������R�ƈ @�l �\ 9���)�ǲ����ߧ�\!�6K�Mil�<���a�d���������_�b,t����݊�����,�qqi�AN��T�:��4RWj�e[�{-c��U#Su�l
�3�߷:���@�]L:u�����_j{|�r��{IIK��K����)�А���4A2zz	e����J|��J+(PJ���w���VΊ�3�ݾ1�*���U=ˋ����~(�S��q�}���E��*��<1Da.f����M��*9e�>}J�ҕ�ș����ޝ�����c��@����ǻd�;�j�?߿NN�*].���Ƚ�%�A�\���m��d�\�k��^�O��&�G+��ׂ������F\��+������<,ƴF�]m9mL��ϝ찺�BW]7^�R�z���L�?��=&~�^�8/-+'׸�j="X���k222ߗ/_R��s�7�d�j=X���0���
����`ؚ��1W�n���nN?!�O�dl�����:�����CV�{R�׊:&\�&͝0]���Ls_�c��ܿ�3��S~5_=;5f}��Q�`����f�\�e��X�v��~���̌a,܅�]�"A���h���Ԕ\Z:��ܥ�h�S��&:۸��\{�noc�7�zC�����e�b_׏����]�#�<�L��]~XO=�a^�W��,�:��>Y	L�՘k�O�����U]j��
V#����n멌$���F�9:�|@���f��`0��������)�C���������~��e���_pkO ���,Q�>��FY>�>e������PI�h�v�u��2o�i����aVG]�a;.�CH��C�cݪ�w������*"	A@5L7�p����b�b˨��F-t3M�f�!�* ��^�	gh���pQ(��&�E5w?�����߯��K<^�4��!0�y�nO@��������x�y��yP�,�>�:�H���L
��Zia�Q��EX]���U]Jѭ�����?��ttt6v�kk��/��Od�ſt�W�B���մIϱ쵱�uO��]5��6¥�������*m�P�g�Դ>��ܧ����r���l�
�J_D��.$�ē]�=�f}W�>��연3o�QTTRRRv��2;�o�),���j��!I�����*��K���lT�^E�Ѻ䫠8�jU��um�|�,�\o��6��O�G�D �e�N旦���o���3=��(*���v�µL�j�x�_�Eʈ�en\"��G��q�������;�T��ml��zǫ׆is�B&��w��s��\f��O6K�����a�i��5UYM�(��sZa/�no�K��<�L��8Jb��l����sE�4��r�Z��#?�,�������4�5z�mvҷD�|�v��S��2���hwӊ~_����LKL��[�3�.����+]���55��>ZL[���}��R�m�5L=�ȳӎ�4�^*D�~Jl�yP`2L���W�����S����D��'3��6Q�2��\��7e��|4����J:#��E�|�^�3��6�����M"�0��6\fc���+V�YZ��c-6�V
n$Y�m����ũ�����2�����)\��l�<�1p��Xu���y*akE a'�;��l�*g�	�8I����o�.�`2�`</g:u^��M���є��+P�C+I�����7��L�:[��A\�;�%u�p3a��O)-�G�5���ا��C�0�V�$������ɏ�l�'�+� �4
�QD�m.���	A�l��e���K�ʺ���2�&��,���`��5l[q���a�\�������/#T�nb��f���kl�&Uܘ����,�f��;""gB_D޽������r�H�F��g���GH��Uk<�!��b����9�4v��-deq�e~sJ�RΚ/+��/�f��?|Χ	�����9-�^|u��5=#���Mu�\p�g���'Z+Q���R�L�?a1>�J�~/�g�^y���?"X�ҝ�.��G7,�5�d��w@.�`�E��-C��)�io�ʜ6"I⇊�b��<�Fr���b:j�O@��m����J%���y||������3�L�F��^�|���i��&����=�Ϳ���J\GM�S�0+g��V?pQ�ig�_���h���;��q80x�h�oX�|kk�q�����Enddd����fz��=��FicxZ����d�>ܲ�kέe�lC�b����� ��'��)���`�	�")����=>N9x�;z�z�]������W�T� �_�i�����������.��yg��^ݟ�'��͉k6 ��C���.,�����J�;7��闓�S��I�,�Nwc�4�4!�>m�Ld�u[�K�J�F,O]�$�
I��3�fQ#W�t���h��N�Rf�e��$I�)�����n|����:�����j�Ը:
g��8ب*p�J�a|+Ek� 34��t����6�ׯ�?]�[=%00���(�_0�����,;/ݳN~�r�H�n+���PI��1�}l��tԇ�������{
��������`��d���ה�����/�`�" _�2666�y��t��N�QBoE������W�Zw
�:�P�?�N*����0�T��Mc�uF:��Jί|h_�9�C����,�D���@�Sҁf?�Ƅ��F�7�Ya>ow�ͼ���y"ui�nt�oal쟭H��~G.���v~��h�����C�N��/	M��7ސy�п�eY�3=&������|�ĳJ,~�"�P�sz�ڇk��6���J��c�N�����:
}VM9���4�r*H�'y��}��_1��b��M�&�Y����~˰��"n}-M��3��T(�3���6���H�٢5�@�C�+*��8o�u���3ɯ>-/�Fi�_^^^t�o�GY�������z�h�^31q�,W�l�e�'b�g٪)�Y�%$Ҕܦ�����+*(¥�_�Nw�Ǿ~���jVp�+�Ib�8}���*�QR�����GE�ŏ��� ���dK4����o�7����3E��WUQ����\ooo�3���{G�����\/v5:&�|Y�]�^*Y���|u����åɠ�ak�����h����������M33��|�N�m�N7=�0�FOfl닳�V}D|��\�%+pqrz�kV�!1��n��=1A�B����¥�܁�~���$Y3;]��Y��C���As�����6�VXb㗜�����ގ��
����X����E����W�u�jY�� ",,,�ڲ������klۄr�%%�k��O�>yF;"@~���_=�� ����q�%\:��_*��o��K��/���ƴ�߿��=�ؙ�z����o�(e�::r��ӟ����)���)))t�Ԉ��Ŕ�\�����35.�>�� �~��t,�u4�ecckL��L,��>ܫE��ױ�H>U5���"� ���[�H���#�]S�@z9���9�p�bM���M�{N���S�\�9������6��ϕ���xs;;�۬����?�����-���-�U���]�g�-�H�#^����>M��C�G3�;�B��៕��E~�ڧl��D�?�����b%�5����<v�k<��5����&&&~��ʞ��vҖr�|�ׯ ӣ4����)��:\�>������ً�9	�~��C��/&&:�}kkk�����ƺ:1�o���OY��7n8�ϗ��~��̈+1v�p��&��S�K���p1��j255��@b��F?�"����#���]> �x��'�Addd8yyo�r��CFԻ���}����Qd�K�����;E���8�H��ޑё���;&�(�s�hA*���я��Ԕ��B�ٱ\[VV6��]��M�%I���+S���9ʁ|���C*aa����z�랞�� r�1:L}�=ql�����v����576h�5\z�9�E*�'
���[���ja`�����gv7�o	A�p9�X���<�h�*m�Y�0�׃�A�h��'g�M`RRd}���"��{;�%Ξ���^��j������JS"������A��bG����RQ!M��6p�cY�i9��^jlL��͛�R!E/� ��2�x��U�F���N��'�[�e����\\��[�{:.1��9Lս���Th�i��XAy�����`u$%�M�7(�[qqq?��>G�m��*pH���'�>U�Rʒ����i�sO!���63��A�ӝ:QB���U�V&,BFA�~mm�Ŵ0���h	�D�ѐ˸�(���M���W�pk�w@����NT��7~��#pp��o��3���	�gY��>zm��	�@���+Y��sq
	Q �;�m.}����n<���o��5��� s4B�>���HB�	��c��Y�VZzp
�O	���a��S_�63A]�q�B��`# �l_�r��C�o�����z�JK��ㅑɕ��Kf⅄׮A�,V�S�2ګ&���[W��t*����)}`8�{�" �����F�aF�˗/<[g�o6���!��	�6z�KN��$�Ȳ�&���Q�D�1g������� $ i���d���襢��ρd��$����N�kjZ��	>��~��G�bv�0�lP���]���0鴲�7� �*�\���oje�qg8���"\XS�'�F����kf�<�i@����._�,@Np0��`�w��U��g+m=5Fȝw+E9:��d�tw���4G���n�z��W�D;�����v<�]z��)�a ��eqL�Es��+�djY���� �Q��>a_lQς�ר���r@s���@�L���B�/u�f��)���M���EIE�"��ׁ+�|�>����%jv��0jp�_c�QUtl�(���ɍ�>�-��(R����j�����$\���A�433�p�kY�)޹Aҋ>#7.X���J����^BT��׃hd���\���ƩF��å �%��X���0���Մ�T�ٶj��'�;����s�oN�H^�oוl0��h8f�@�=::����m����ίi2jj����I���砓��Q�},&H��*��Tȷ�J�SCh��oI����] R�ӽ�u��WA�.G������9�f3v%��{Q��q�	b|�����>��n�K~-�U�r6H�)�L<�� �
���w�@�iθ�y���[�g�^�'>���`��[+(�{੕v-��@&9���� �·J��bnc��5�.7�~$���4��sb'GO�*k� ��_~����5BAP�7q�s�'��#��{�>������mB���*�4.*���Ċ�_��7[
H�<v��k�_��B>~������`;$�M����u��R���UmYY���`����Q@ �;�3Ȕ1W$�����N�����޴&���~�@�99��; ��uƿ����E|��i�<���׿����z�Z0��� �Č�t����͙
���^t
?��p|�X>i��x��ѕ��0(�l���i�TV|�5���c��>C�]��dR!<�
�A꺺�gI��v�4;tk>"YFs�҂�~���wڹ�����1�a<�D�	��\�̪*����_K1㕃e��}It������r�>��w:4�����Q�K� ��]�FVnW`Yly���f����;��\�?�J������.��7���OЀ?�~�O����G��N*Y٢T֠���W��B��P�[���OБz�����M�� Xp{ХN[�꪿��k�x�Ĝ<<7+]0�?��s57�ΟP�y����*i���GS���D<��:`%	��QRZ�$�qL��!�p��;���u���]�(d�F����:g��ěPut�!2�&��3�n@�N�=�{��.�������l�b�I&)���m�sr���P8�$ZYY$����!O
�H�(@y M��g�V��F%�G�a��,;I#�C�bN7SeDó�vbp�U/������I��w��V��"Em-��K� �G����L�ݴ��b�?������\Q<�7��-���m]8.	�⯧�|�p��K{_����\Z\���R��V�Ύ+�G�j�cS	�����)8�<��9��6{6ZB�+"_F���m[��ek�n+e����'�����һ�J��X�c�j�� b�Eƿ��V�� ��0�}q@�$ص)G��3pu��ǧx�!q���A^>)j���pv����O���l3֣�� �JtE�4�y!7ܹH�~-��?�B��yu@LN�!yz�Z��;�cV�����:F���P�t�u�IO�r�{�����B��g٪�^����*}�Vc.�_S�-󎄢+___��!(~�Z���;�94S��'>�K��O@(�C�����'�/@N6ttȾ�`]T$>>:��j� �j
@��KU���=��p����`�g�p,h]6H�t6����6:@W���$~����^\�8���+\X\���S؊F
a����T��]��4Ֆ��gA��LZ����ozz��8zcdX)��/ � `[�E���P�qP]�իW���ssr����M���~�4m6a�4���Q�~i'�t�uB �Y z���]� l�Yk�X�ѣ��s5�����ٙf����3`v#�?8�j�z{{����.��
e�  @�y�f�=�3��N�e���A �y���y(��.���?o���0d����M󽏏�6:� ��nYL�W ���`� ���XX�0��pV(�>;f��"�pI��{�w�#(����t������HB�Q�e����?H������p����l@�qm�0���<y23V�BN�T3�	� f��H�7��р��0]9"I��(�Z���������\iU�A�3S�| 6��!�%�0Hb@$LVʔ(����xzoYm��B��A����# ������v�*{��#�Ė���+�K��JV?�<T��4p��]'��!d������ jM	�3 �E�>��#�Q�5?=���}���uǳ3_$�1�Ùå9��9����o8���rx��$-��05�mK#�0"2��As�݊�5��e �L�q�~= v�N�=����e*}IYY� #=0W vH	�����oZ�Z��	�g�UB�-WX� 2s++8�T4H�oD���O\�1�vzR� �1�/������-.)�P��Tw�"6P�\X�}֕3�+כ)))������h`~'~�شB�"�j<HuE�>	���5����@|�m���������/��_�����D���x�� 9Ъ�??�=e�zNNNh�Pu���/㢑}8�&?d�)8FN�qW����x�"��&?<<<F}���LI�G����� �Ƚ	N�X{��1
�|#�T�=AN.u���q8���(e���� �I����ߎ��
���'�Gh��l4�8�;u����Up�'�H��9D��?��@���O��!�����;�2��P���A��Q>��5�s]*R!�����@ �{�2,B6���V������d ] ?��}>���j�nR�9��ܓ4��|�'Tq7�UB2�m!���v�D5b���^���w�lq�����~U7�G1E����jMa��S��wf��JU�k�M����
T�:Ju��V�e.���?g�\<�D��E���,RhXNL��H�@5��������dX��o�?�|>;��oƚe���>Ig�Y-����$%L����oG�kC�4����h�o)�]J�kw�.�P������Z�D��BK��"�IgC�bN���Q5�4R�(,�֊z-�b޹x�W;x-(�XĘN֩,FV��=�#�`h�^n���1׺K���6�m�=�[�LpU��ƷE����o [_���%#��}Z����x&��֯O[����]�/f���tI�Gc�3q��ލ�؉��M��Q;ݤ�|5������~|�cG�:�k+zǯ��5ۗ;-j�R��-��i�_��NArzeu��s0��{hҪ}~��s�����#�eI/���L����+�)W{C�x�D�&����VOG��z�h�����	m��ե �%b�����z��$�3�u�1��0�DC�}@-z{0��m�[��O�تt��>��������]�x�P=�����Q�i �z7rT���9�7�%��w���R����yRk������u1����~��T�x�`����� 1��ÆB HVaI;��c�e�붱1�t(��Ӧ���������\���%/�7��[�������b����=�[Y^~���P�8��QBO���ڃn��XĊ�~.��tŸ+�oY����6s�moo��=��=v��8 ��� d���\U饔�[��������$6�ik�gf/�v���
�Z����������˱\{s�6ۅ6d	-`�gf�������+Ǔ�u�\�O�F5�v]�ܪ�r@��������y��t"Da�\��=]j�p�@��5nr�*l��@bt�p�(��?��C=�ֽ���{[�E����N���G����j�)S�>�^��K&�d�W�"Iff]�_��`kЗ�+�_4�f(e7ez�9:کm���T�������{�e!%����}s �o���\���Sz���B�f&=�bf�kw�@��?vЪ���%��M��A�Ӏ����*���At�q����j;�g��E=o����E۟F��kׂ]��h����An(I�����@����o؇����%�klH;;�&�Fڣ����tnlH@|��2UΒD"�z��C;����'ڟ�%B�vk��r�����q_֬�Ȏ� U�h_�ՌY6�n���@n��hv��7��M�p/���H͐*������$�0�C{�JM�j�M�����_��m�+�Θ6K�����5�ބj��HR�>ĞaՁ����5�a��h�0W#�F�v�FG)��9���`rz�U�m�&D$��s(���[�q�$f�|y�(.)�e�+l�*����c����ît�ÞKGHL��z4f�~ѻ!������srv~�#'��%dk9���j�!{�~�����u�[n�?:W��r��� o�	�n��c�'����ǈ��
w�l����|����	@�ѐ!��KU=�}����uϯ]Ci�ny#7��h$X3����hVcv搳�	RᡠjL���L���L)�ܞ���� ����8���>d�Y_����C]x>{���h�6�Z�`7�M1G�6�L�y���S	G{�h,t�)4u���!�TSS����ǂ "0�2+,��i�T�7�5���7�)�+���*�L��F����l�ˁ����6�'f�V�8�)���$4L];�e�n��-� 0>8�9���K�z!�eu�}���H����q͹�A�R��Eg�)��Uq~��7�}'S����OL,q�1.����i��qV��#��/jl��3�J8~��=͸�����J��ᗤ[[��X�u@��5�o����m���}W��H/�1�/�5�ޫ�ܴ��.q4���:T�u����,�xQ����}����d�O ޥ���.k�w$�z���<G@G�L4Z�%���� 
'�>O���%
�GYK�˚��_?Oo��1��I��V�"��Pf��~�^�ڞ�^���є�7�Y_�'�c����\j��&��җ�E��e}~̿�=��{��%���D)�������&T��C8)�P�n�<�HL��X[�=�k�K"r @߀iJl�v�mq���<Q��e����?�A
���j��s�[Y*Y˲�A"��g�IR?Ǒ�>��8��8l8�)a�i��,fx�@PtR �Low�����M��Cl���+��I������Y�!� �JZ�|E.�c�/���N�1j���va3�J|+57�2ߞc3���ز�q�%�}pv���7��j��Z|k�fM�������c+�c�;;[���RO��b�,� <[���	�L��Ų�����mD*<�p�c����+�ȑT�s�H�R� z��s��������𮂊�����B�͊-w�G[�Q���B�#~����IVSI{����͓h�A
|/[�������s�'o�&��vm�{��E��F)�7~֠[;���+�:�-���&���t4?�lk��p��`M�L��~~2�&���̖k� ��qC4�<�Ѭ�n����V��p;!�f�6���_���=k�	IIIHR�~'%�<��5F*?^����b�����ir�{d���q	ѱ�%�)�B�^f��W�`w71v0
\M�c�s� �1Ķ���-Q��0�hrrSX���'�E����qU��SF�D�+Y�_���'�b���{�h��$�jƊ����&��1;7�	�#�@�-Dc��oK&zG��
��PS� C2�����4�ʍ��D�K�VG��OCR��=F�N^��`�B-���B��������8�X+0,333 j��������S֌��?�����
O��4:n�M�Zl)!q��3��N�&�<���]�f��4iM:z�v�׏�h-]���^��z��Q�N(f'��t�h���NK�D���XS��}m��T����.�|�nm���j}*�II�1��Z=+�1��5�_/�����"��-�b��v������M��$������jX��.
���o}���m�CLc�<�V=�u`:�ںjs*0n��GO=��Gg;Zo�L(/mD��q�k�ۥo��	Ōn��(�r���ʽ����7�{��碳��?�9�ϥ�Pz�6�8��������#�:d�'���T-�)�*DU�P�̱�<GAO�f�.=콟9����s��լvwA�H���6�Xu]��6�F�J� :�(r3�rk�y�w|����I/��me��f��s����C��9���#Z�IL���I�;��r1Mj�� ����8X^�N�ޱ(Km����}��P�n)��mz�sV��w���U��y�Sa��Ϣ?׮���,9���-�/���t��S�VYe[�Ń�:g�{�cQH��R�����C�m�3�ۥe���KL&{>��(��q�픪s�;��U��n�Ţ8	�tk	6��of��{?����h-��؊���j��QMp��g@W�K����	�p�e�E�
ͽ1zz)G�v�$5�'��� ��-��d�,%��?�m�D�D^&�s�e n�iZ�˂��x���I�(��;QsD2)�Yq��ͭ���'�
�D��|�~�h[���kL.`�`��uf��}���}?k=�2�ܦ׍�'mєG2G��
s�Ǜ�R�=���<Q&=/�۹7WE���^���&
��ri�ݯ$Bq(^�����F������*���l2�[j��Iy�|	�bU|��q�E%ܢ�9IS�
k� ��$�r��<w��������8"Mm<~c�b����Xg{m�Y�����z�H�I�Q��G���f���	��³w3���iIH�xm��y���伂
�W�?(i���G^Q�d���+�}��P��>�*G�O���[\��~)J@#­�������(}$Ad���U���&W�tQ�]��G3���}�������z@TB����",���6�`��Tj�L���笄I99�.E���y6z<�8���^�q�#>��[�9"4���0'�óck��l����b)rB/%�}�L]wF7�F�9�QL=�����_p�tn:�ˬ��S��`L������]y����>����YWA�q��lS	)�u�o%YFqy��Lz5+�I��_�	��9��&7l��!V��6#��7.�b<W$�U�����M�o߿��`�<U+���/����h���H�QeV�h�[��������!�A�s)�>Z�
?��j��t�d�XzC^|��[]Ʒ��Z��3~j�lx�s�\��۝֠m���Pf�E�c���\�c�QP��`���.����K#�x�5���%� j\)�z��U����a��:��i��H9݄���g�sH����:q	�5�7���3�����{��*#�gG4`�� N�XS��
dZ�gy��Mu�U����VH�i�2��̍����"�m�dnv�����
�qp�<�D#��g聈Kb��:�	8��?=Ikilt���ȹ���6������Ԡ9�	Jm���HDy�W�R,HB���0~��r���,UAe͡O,n=���#��*wv��ԏ'{��t�b���z���3E{c8H�@��N<ჸ��=���x;nPZ���u�����J5�TI�I��p�aT6�i��¹��Y����O��֣"�{}[�}�>I ���A >�j0��2ģʢHE����bn�h��0���3Z���]�y{n`�[[�X3J���������ZK�[yp�S8��W���c�!�d���ݶSO<��*N X�Y^���i݅���
q�B݇�d9#�"�I�d��Q�u�d�j����Z�v�#�nQ�b�Ŭ�U���	��_�	��/����4������`�}��/v�,�]T�ik�nJ�#��+�ƋJ��H�>��Ӕo�Sέ���=~��O�p�H0��ll�8���u���G�W�2��&���u&k�Jh6�C��v/��������y��:j�?~�ϵ70�qw�j��_̎� s�Z�a!����c{�6��h��\�'i"^�5��˜�
�^�do��"m�1�^z�ax���a:4A���7G�O{o��|0��G"X�����X� ��+$:2-?d�[j�+4���n�Dy`��_1z�-ҺTx��c[ݔ�C�y^}��#��r��9��9��l�[���o\:�����v+�y��KE ������]LQ��Bּx ]Z�l��9�; �1E���&P��H�;`E����o�&�#�ݜ,�������c�l�W��|��}�I�e�6B{=����Hf�$��&��휘w���#�Hi{Eun���ư�^t�(��԰���KK�k�԰��C��^c�5h�ݛ^G/?�(�#洿�蔡��*��5P��`$c�[-m�۶!�y�\"�����X��>p��%h�#譞L,f�]���`���^u����������j���]�%U��!����sƔZ#��^��7UZJ�u��L4�p��T�b�]�SO�pcU�[���L!`�@����QZ����Z9*���uX2��]���o/��E�Cw��L�����>�{�:��R�@:��E�`i>GXIʆ�Ҙ��`�o��+�4:Ô�_3�5g���?u��������й��E~�s,���hN��+��8�j�7b�y\}����r�5+�%�T�O;���RA.�#�����B*l���S,�w ����X�wy+0c�#5T�C�m��ƾc���Aa伄�|�������g�º���Rp@$��������/�Dϭ2`u�3Q�a�+�<l�.�x����������=�IÈ�J]?åG믧g�}7���]+�=l��_�x�>��{zd|�����+��+��g=��F\V2q�Λ��@�6v*��+���Q����z~0�i��)잁��m=�&)��)�X�������^C�g���n|@��\OvϯG�]�r��Xh��a�D9������=��hhj'�E��^�3��pMІuRr�@�UxB�æ(�COɘ=c�A�s����"�"��k��y&��wv�6�8_+�?���ߡa�	�Ez�� q%}�&)�ӧ_���!*�(~�xh݊��47�<闁�ϟS����p����*����	ˆW���S���ёm�}0�w�\X��V�|�gM�+)6T'\�p��)���������a�O!�d����tS7� mT|~��#z0B�@|�+��<{����O>��Ͻ
7u�
�}k��#�U�n�v�/�7Of��:̕Zo��f�b�}�������P��Z�䝒�]{k4���`IA�� ��z>R���};��[B�7�aN�IA\�j~j:�(Ց�jJ�n:��v�CC�	+�Q��76�Z8��&$]Q8���z ݑ~mˤg?$��{z(�'j�o��Nmd�5>y8�B���-��"-ک�'�m�2v�����ؼGh��/�_�W�"Q0܉�=����@c�P�?�9�74=��SO��f�����]�L�ޣ����@"�V���1�J:���+?0/��8�/�[�ܧ�O{o�{5�^����O���$(���8��\2cxu������yQ��$��2��
-!�#A�^�)�S�������sǭU�4���xd����G[R�RUp��O���+/��6��;���u��|q(�MYE�GpC�qP�Q��9J�U�;<�02��J�TU��#�ǘ\�L�}�dqȿ��	�Ȋ)�V�y*)t�A>#�F#O�4��a۱5[e�[:moǽ���|){�@�w��i.fgZ�;/�^w|K*���.�:���8γ�RI�]�����w������.��{��Y_H�:��[�*�%~�(vy�=��2�u��j�e���-^!��Z��%��6���{�����u'e2�F�F���Ā� K�sݮmIk�ˊ[sa���k�p��*�6�m�t	����8؉���h����T3��mc��|�g԰u�$p7�9�n���)���S_n��ʱȅ*�����'4t��:����ò5�#K �����
�JPԴe�x�Y�����؀��r
�*Ļ>���˹�--�����5�\{�f��Q1յ�\�I��Z���}v�5����D����K�&V���+]B'����m�Q��1�B�\�;�A���_���,P�7�'�!�q�`L^��`��a�ZE��U;BNU�`��ff'���S�{�FC��{3�tWbl��Vx�Y��^����x�'-d����@���R]���5%5,�a�Q�}�la=��ۓ��w��Ze�<B	4��7��L����'�ٱ�%��퇵�|��Y�c`����uq��~:R9?܂{7�:[7�;b�{�9Ɵ�L���\1Tx
"m��v�u"'��zޫ� �.4�����z@p�s��;uA�;���
4�>����N��������׺��qs���7��BNb�n��j�sI�����?�e�xX0dL��5�ͻB"6͵�m၊M_m�jU��^��&
zж3*C���j�k�u���_N�M<{>Xf����ͱ@�*$�������ɬ�Z�X�k_�z�]�����5]y�+IUi�:D�K�=
R�'���h�O7>��+����/���sU��
����1�W�^�U�7hg���_�J,YBo�Dd������!��mX17��MuDW�.�O�S�/�����?{Cv����*�s��m��4��?���fZ"���N3�2�:G����+!����2v7�8��J���>	��%�g��B�^i�\�~��fŸqo�o����gW�ɽ��j�ωt.�-\~��V�[FyѶ��ho��N�k�[�o���I�<7V�B=��v�	G�v����_�o����S�!�_y��U��� ����S2r�b;���W�M;�_ˌLn��C&�IW��mw&Z��ϵ��4�C=�!��J�\��E���C���Mo����p>�}p����'���7��BD�:��Z�������2����{3��hܩ�GM�fX?�s�R�%]Be��߷��kr��"�Ll��GNVz��Xk��N=.�4���'�rh]�\)V#�Y��k�����\��[/�l����$�7��>]	%/�ڊ�e�jg7����N�4��\3<���]C� GM��<�ͯUe�D:��Z�����&I8��%[nUm�ƿ߫��f*H2K�{�8$SK�ߪ������?:i���^�W��b�j�e�qd%�鞵�H���~	�C׷c����M��v���x�A"[K�Z������ɽ��R��u�T�Ӟb��J��*�μf��k!a�}�M˻��S������p���vF�n��J�[�5�����>����!�VOO�D�֮���Qm��6]�����Zd�.QpJw�����$v-���F��ˎ�\r��t�7{�zZ��z^*�R|�ט2:��5��9vd�N�z�>�Sm�3תt�	W�Aٿ�7��Y�6�0F8����Vk	�����O�DH���]���7��1�������.�A������+2���*�7�P��ގO�ꜚ�h�Y�ֵS���F���<Q`sO�`n�-�I����/��V˨�?���z��?��s�X��A':�/�Zk@�U�Zߣ`YZ֝��e�7��[�U��,��JI1�{�9�Q��)�^����Sn�펍���$��/A	��L�w6	ɬ��Xx`+Z�Ǯ�ޘ��`_�͐>�q�?��^��P���S��!��C�K���&�$�薊��=���WH�4��8O-QZ�H��,��z���^c}�C;T���󊫈?ܷ�f��V���#*B)U�52�c���1�g�-��g5>�7?����{�tt�^(�;�1�%�1���鐷�Zҍ�~��H����:#H���GGu�Ũ�����E�~�MU��{`���63�Ar{���n���n�z>^��v�^���)����	<�a���ݑ�q����ž���~�L�;�Ą�`r'�hHw`�v�C��]�yiXtxi�����s4$o���V�������Ki���V�VǶ�.S�w��Z�e��.��`j��g�I0�$a�o�NV}w<\g�-my#<R���r��~̀�����j�4�w��UlS�oWL�J��&?���\`x8�g^���t��r�⤜!������j%��h�@w2(�F�J�9��MSV[/5���5Q����A���9��������[��UH��zZ��1���Ⱥ�&����DiOi�ҥ�bA��ҋ��� `�J�EiB��@��ޤFB�bH�	%����S?��x8�ν3w�73ww��u �zǱ�1D�Y�N�Us)��`�m��=v�����[n���"���&?-j��Vh��	�*�<W~�<��?\�4�@��X�W}��r*���F�S�������%LYr� �f�ȸ�3L������.��2��	1揍�������e��Q�.�����)�m���qhӾ��y��fV���*cm?�����$p���8ʩ��n�i�o(�5M#{'�0I�T���#Jo����U�������(�z^nPY�L����Du��[�a|�?�:ĳ�,��r�$=X˝�6֖�p�mT�ɟ�S$J5J�P���ޜ��ѩ��4��cL2�P���q�[�s����h�>c��r	����������#��������UW�+V��;�"�M(�7�<�1���X�|p&O�c꽼��a��������/����,�Nmۉc���R����F��	�_#'�m�Q��yѺ����;KM�����W^vtɎ�H�9���"����Џ���{A3P7�}�W�R=���H�/�c�ޏ��vp�1N�G��yW��ۚ� #�E�Հ.�kS��'<�#ɋ��L%�~��t u�)��>4[��賿&��$e��#�v��`���&1]X_�e�;ѫ� �S���.=�>�ZɳLV)���z�!��<+l���t��|)d�)]mՐ�
s����m�`�u&\�j�q��3�R}��;��ѧ#�D�#�2���j�cA&�}���i	j�14h�}{�|�Y�0d�	?,���G5Mnƒǒ�M���\3|�Q��X������ܙ�?.����MY�|; �� �o?�;E���$��ќ$�}�0$WS������'��H����e�޲2������5���q���)�ma�x����8x�E,�A�/�a�"�����V�"l��B��L�'�P��p]�U:�GI/���N�U�`���x�-'�Ӻh���GGz~�=X�a}�J���� ��аo0�O/@�*P\1=��pu����}�i�: eӺY�{;�����@��V�H��&oK�MY�9巂󬒻�O���A���骉,k��x/I^R�������i�L��m,�g�;���&��B*!�
	-ͦF���ը�x+I���	 2��-b����4�U�ᄹY8�l��&��Ĭ��?ulw�p�f�Z`-�(	��|���Sq��!+y. ��rt`$i���$��JG,'���p�1\�~��cIY�����&��G�^~5!z(������7��8�&�88؝��,p>�p���CV����ek��Ks��$�mH�m�@���!� ��:px�MBl�{�Ա)[���׶T�=�񟉝/Y'K?��� #����U�f^,�d>���+���f��V�1�����U��B�����4����)���z+|��x��crN�����"�'�������i�T��_�7��������!���W���������ݞv�5�r�Oώ&k�g�Mp��Լ��)$�-��f�d�=����{_��$t��5�̬�w�e(�k)������I#�����]w�,����.]1� }8Pn�B���#�;��
4BpM���=��C( A��A�>���� �)#Q6w�Ք��O�H��,����Z�Her�ʈM��GS��� ��&��y�8K�>�����glu]�Nc�1�י�TGk��V�DD��wPIL�%�G���p3;/IRj�cIxu�*��iu}���k@����8��B�����K	K������dZ�"]ԕF�L�>ߥP�����gc��@Ѷuha��?8O~�_W�<��,k���J
�o��������̊n��T�ɛQu�̸Ք�����6��Jd��=D����R1���~��H�����C9$-W-P�J��B�D���V�B��4_�I�Y,�e����_I�`�I�}�|K�7?3�藄0g�����KQZ��Ő�~���� ��z�E�%\-���_60S�4A\����zwf�\�wA.]�-��:Ghnڎ�36��#	�=��{�w���� Y��:O��;��sjӓ�чr�B��=đ��K��7�AU��Eoi�,��{,:�4�_��
O��.��i�s����	b��Ey��M�?),ˏ�h}�^M�v|�s�;y$G���,���-����1��c6@"�6r3���f"_p�=�n����C~3�v����?��m�_O֮jrsS.Tm���Av�j{�< ����M�^�3[�9hi���Kn�Є����#��"�L#��I�nmE��};wϻu7�v1'ϵ|B}�L�e���m����ȯRg�2,��&�Wƺ��͟����[d�A��	�9 Td�F=4����j�:��ma��߳%1����ܐ`յ���
�,���9`��pm��>�DW�I�Dо�V� X:��O�GɁ����������e*�:�&�A,Ca>f�\fKJ}�w�~%��8��\@�W��U��$�U]c���_Yۀ�N�̅X��x6eU d��*��A�T��ٟ�W��Y�\5x�Gn&j�S��p̶p�1I�O.�]y��L��]� O�z�<�X���<�|�� _�*�� �F?�y���5��F�6�LM ��=�����~�Ќb�!�_g3���n,>�D~���(�J7)�zz��q*��q�fTkV/�z��k	��q�TfY�k�j�]!>������3���;��_�("�4 ��{|�j�x\�eQF0"l�z��Q�M9oJt�����RM���F�j�\��]�Pf{q�rS�e�ͥ�:�w�\ߪ��u�Ў#*��
��iċ�:�й�k��'h*�� m3�E�~k����
��W35�v&��ՠ��tS��5xuY
��LB��s;W��~r�bsn�*��	��)�u򚒪]����Ɵ40<={��2w���D�Dи�r�a j� �b����9Bl�
B�N� ��Vz0���D�O���J�-d�-nz���z�C�/3�b}��},F�{](�m�ȍr�͠��&$=��]���1o"�C(��μ.��	c�/r�ǚg����yVY-�9�Ǝ���5]6�|.��	�]���^�LqAq_��LW�ӹ?�=�V׶�q�o[��MUE�SV(ࡩ梪ôcxwqKȒ��D!r�7��n΢�Xݛn\ǖx�b Lo� �ޒ��]^���t��������Q��T%����߂LU-q_��2�����z�<�V���R8k]�J7 ��8i����ΡN㱚Bgc�ܻq��߿��癟�x0P��p*������5rn��c���J�����5Q. @ ���f�6����3^��<�hBR��d0�Z�#���et������]���G���DA���qn�6����{�!��ަ�(��n6��q�^D��B,KꂡC���ԬQWv��`1��a��'�!�ِZÎ׿���aj�3��]���r 3�7�>xo��k�U��#���s[���D�\�	�QK���~��t�P^i����d����:a��.Y�]đ�6�h'T�����߂�#������$�I6���xs/��O��7��@W�WR�{=�@�2��lz�� !��}Z��q��Q�#V-)���D倨��!���$�sȹl){�$fw?����� ^} O��䫁���ī(ҕ�0˙��ܧq�I1�Ǵ!���2lLU�h�qI�v���v�T/�=�]V�I*�,�X m�k��'����F�tƠ˝ӣ�B�Y�8�)�^����l��Lm����U���� �ء��B�dZ`L��*�g֘�Y�BK����e�C�:�+�e2W��
��-R�&<.)Y�	��Ȫ��A���DP՟H�:�52<Z�0xm$n��W�\���������G��l	�UVN|l�E(��9`�����Cg�H�d��.'7�<J7R|o����+g�~�*���ׂ�-��e9ЬJH�b��R�!��Ǔ�I2�^�C��RK�o��b�蜚��=��gј~@��y�_qg�
d���|Yl�9����z���n�՝qݧ� ��ӷ�1̜�v滝А�YJ�P_�	'ip��G�o�qo�P��蚶:��{#M1Կd/�uG6�}��fQ�����J&�_����rD��%��"d�f�ӣo^,���7�i!}��h���_��F�Rԃ&�V��[�M���nt#���yLfе�d1㖃/�[;�(/0(e
D��|�Fv��V�o�����l���U_൴kq��zF�Z���� ׎C�	ږ����Y��ü�]:�a���[� =��|\���.���'8�mm�h�U���y��`P�Z�{^������6�����;�:H����濪/$J)�+��Hsđ��+��=��3�|^]>:ﵪs�A��7Ϩ~�����N��a�H\U�A;���8�͕��������щ�/X_�j����ٔ:���oNi��A�@��gmt7��"P4���.�jtU�/I��~��+�{_/��K��4]�}e��~��X`���2�o�Q}'$���48��ax��Q8��^ƞt�Vn�50�[@����]U�џz�/���͂{��TB�͹Ǡ��.W�]AZ�8��p�ąLJU���9r�.�r�ii(j��7@'�(��T ��]�2���ǿ'AG�ٺ��Tp�H-Б+̵��呕լ/ͫ9��$��rĆʒjPx��q���Q-���ݹ����]�#�����JK-���x��:���~�OW�e����E�!��NFN��A>�Gm�)I�S����.�zhK}.�ud�j}��گ�����s���1O�1-M�٨#��_f�)c&~���,�ϧ���A�*4b�V�@H�ĩ��@(.katW2q/B��˯�M\�I4z�T�4j6�6.�=��a��!e#X�3����0-�N�~�P�_�D���i��7�^aS���>�R��I��o��JZա��~1K'�o��.}Q���n0W�ee����z�yw��U�<l����SC��#0���j{��ݼ�Z���q�~O��^7����5���t�}5�b��c�@%��uy�4�}�h�o�1���90j��!hc���J8�2���ї��W�Es��G��s�P�xG�[J�U9�Ү�H�'
V^�2�q[�U�l��h4{����$pp2��D;WK�4�J��m>9�~��/�V��XE��7C�hk,S*�M�z�]A%�4�����^�f�1[�}F7���ȇ��}����}�?�}d�s��~���{p�Q�q�-�}�z�AveВ�4�#| ��ӽ�}�o.�ұN�s��Śf�
�O��Vi���Tl�����:q��tS�;�ٔAsa��o�; ;�q�^ �4�h�����9���;5�A�~�$׆���Q@��:bs��Y���ׯW��w�b�-<���������>����<��r���"w�oCx����y���<�2��`�$;	hk���L���:�q���*8��p�LlLo�@�A�8����Ep�Zpl�a����!�A,�]#�Am�ă`C�����='�w��x��8�yZC˜���;L��p��~�1&o����)ov��������0/�<��NB�pQE<V4Ѷj�~m�m�=#�!���h�{��E�2"���A�<n�KW��9�5<��'�ǻQ\M��l���o	��T�ȥ�WiV@��>�?�rT�	�ZP��C2�|�����5�����i�����F)z��V�X��RU�\�tCS��5����\�1&�~e\�d||cF�n�ͻ��)�d�����b8�u�&�n ����5�Ԟ�Q�e�X�!o��$%�ѥ�w�ޑm��Ȍp�����쬓�S�ɸ���||�h�ag���	�v�^N纭�2 ��Q6�令��+l����M��]�v>9�fxz�نChN����\<���?�!0s�z�o��P��L�Ɗ��#���j�9l-���/����)����F_���n߹1���\���i�>s,�ܝ����2̾PFZ��VH�x�8�xT��'2��0�C��Pބ�Y�U���/Or:o�X�����EY����+l��n�~f��I��R�K~yA�Q�(_�֩�h�@���qoCW���i�� kw�K��� 4���O׋Kt���9kO
xo��W(�'2s'q����P��iO<�0R���*E}�WL�e�k;����s�||�uܿ{&A7���.��9O��4��%i<0��
���m������[��a襸j%�K�1��Q�>�PYhcU����ԡ�J!��uW�e7�W�0�;�LՁu��6d�&|i�[�	c�ǌ������x���8>[��]���GkƯw7�c�j+	}f_v6�̯��@�g�_پ�*���V	�� LE��{^�Y�5��Ƴ��mt���^e�Uu�4o����;:�QpÅ������g1�՘4ʢ�ȩ�ҏ�H��m���ҢsT�`ĩ��6�I&�3��+X�l	A�,Hۍ&f���o�Y¯p[�=$E��;����q1��*��Y��3ͻï̝��uF3�'7F+���@O�"�o��;�PsR��ٯ�.�5�:�;`�jq��O�f�\��3A�5R�n���|ś4���g�}`��wZ�.Mɘ�u����*0�pJ�En<����`�o��6��p������SZ8���Zh����8Vo�QXm���:��o)�}�siTB/�K���������Lo�U�\ǎ+�1ѧ��/fM�suo���C�y�Z�)%�}
�fk���WKc���y@�A���m��m���W9[��]}���|R�cuv��ިx5H`��,�|�����h9&\�O4�?��d�/c�,vR�ޫgr��m�����t���a�?{Cꐎw5p�h�+��$Qt�6��1����^PXX�u#=��nx�� �H�)]�O�|�91�J��˗J���U���]�e�?�8X���=��X~��ʮ��F�������������m�XnI�n!,m���Śk8ƺ{��%N�3��7��N�N!��7q�&o�	���6��>%U�����c��gQnh{(�֑�s�aw��q�Xix4��i�{۱����3��_#J.r�N�J��ￒ5wK/^q�ZV<q�A���1��4F��w�xY��I��zy ���n~~�b8�nJl[��k�H�W�[NA��erd+7Q�������4K�n�/=�xV�3mV��Qq�}������
�73��%Ť�ry`J�&������5��S7q���e
��2n�fyN8�4�8x77��ѡ�w�
�6"����|�zR�ⵏ�<�s�+�Q��^�����'|���隵�?X�o&|���YX&��x긃(�<��� ���a���VC}�S{�Ii�yߵ�M�]"J����^�u�v?EA��T��\�$�n����:;���wO���ox\f� p�ڄ��U����e�Ԃx�m���?l����������>���o!�z�R�q�0�T��aUqT�:+N�uQ�f�t�݁��u�Y>=��A�`�]�պ�:#��Ǻw��&�b���RH��0�_�)���q4�1���p ]�}nRޥj>�[��x�K:D�u ��F�H����+\O�!:?�[ȼ�a������J�u�P�Q~�Cc؈�ѱ��gBN���Y)�ڡ.6��QC�UU�V�����i�r�5��{`�!ڌ%����*�������|��v�h��1�͌	�a����`�'٥jF�z�8����g�ui��,���xx��nz/ؠ��Lܰn_�g4��)%X��e�	#��"�Fju#��ŵ���y�]&"������Y��� �r����y��Z�##h�$qss:c�]r�C�f��vMtZj=��Tc4�gxߦO�]9��Yyq�����JI�踡�����&S��mOii	��S[j�Cr��ؠ�Z٦�����b����J��'� �/��>&RD\Fla��R7��O��N�w阰&¦ �3����$�SL1��S��Ix�����q�É|�ˢ��r���n��e��/��XY��/��!�7�jxI[2���a}����)��^{�5�XE�81b��c@y��/�T�s�"[�CI��_�<+
��0�O��&�t��615�d<QF:��md�������p��c�~�3�~u�{yp�u��7��B����]N����H\�n��_���P�}�piBx�8f1�BT'^ac��^Y��i��/(�N��1�1S8�f��vq2�t�S0��2Tx�p�x��R|f9T� {O]Ҭ�m7X���G��;7����v��KJ��
h��\\_!>�b1Oҽ���ZX��6F#�GT�wc�u�ܸ������f�)2|�[�PȞ���_��6����}����c�Io��_ �AI���i�]��&��U��jB�%^�z9��{���m[	Q���h�j/E�2maS��h��F#F�)�.[�qjrg��嶐ܷ,.�K�J�h�8j@�OMz�S�������GC�����.��كc� nP�Fĕ� ��p��'��1M���w��U2�wMK�:g�I��8݇���ǣ�{��}�����*�kX� �s�;=.���|w󣫱ǚ9���R2����!�*�&r�y2���i��
�M.=�D�-+�%u�M�M����k D�O�-��k��"Uʫ��Xp�`�u���ʸ =�q��U-����B�� �Q��\����^������lE|�
b�n ��Ӱ�Jڛ��9�h�Ӑ<�l[��b��k35+6��i�I
����X����G3o��(½q�=��}��s)N9����ު���:}�=��2g���ׯs���ְ��rVoXXح"���垟G�4� ��F��Ep(T�~Q{<�,{@wR��%UA���2n6� ��2FD�n9nw�)��7�,uJb�U�b����ä��"�j�0ʉ��l��v]n�������dgz{i��\�ç�T6�3�v��ґ6�;vT�U�o��_ hD/;m��j��?��^JyV��Wi���*q���Q���j`�g����c�
�Vk9�kv�������Jd����P7l�3���x�놐;�մ�x9B3�"�U���j��ˈ�-&� KOlrҰ���A��T�s��y�<PuϱT��"�櫾;z$ʁ�'�;(��h�Lo��b��#��S��t�U��%a[Y�\�2�A�j�����6-t �vr	9��D�#έJ78��R���܎9���0�K�����f�s�C�J�ѵ�CR-���:�iG�mmn��v*#�7�9��FB95�ћ��př��뵙�K˚8��2�0��չ.*��]elɏ��\x��b��#�%�B�fr+Zg�q�����o���iY�	�!4��z![��§�xL̸ωn��2�%1��2'9�t�,��!�&�I4��7��\������k���EC��qP�]�M\	xǆ"�ګhs_c�1:��X���L�.˗�T����W�ȝt6q�R�So��#�8;m���汑D��g�����Eok�l�m~KS�N�q[xr�f�k�".�cm�;ó5.$������������m��3��d�Dh�TL�?���|�W�d��%���5���8}Fs�mL��@k����O�ҾoW���(�ʵWa`m�;��e
�ћ�{����i�6�p�P�����q{?�/�y�U��f�xgў��O�LD��A�j�M���:U���+�PUIc��8������#�!R΂��cN$S%����M��Did�V��8:����ns�R�xĳ�AT1m?�)x�+�^�C�z��ǡPwh��ǅ���F�9��{?��~�!�d�U�����)��6��p��A�@w�k��u�z�T'J.����k��W;�<�y�]�6�+���~M*/O��|��m��π�����\�2Co�h���:9k!��;�I�V���ou�Q{Sq��|���۰�4pȀ Ug����y)bR�j�:הQ<E�|f2���d7À�z5��Z�a�k��| 7���!���&yN���^��?�t�5}@�ԋ�X�~��"K%���eܧ����2K�Ճ����-�4��0iRxru5��dS^��y����2mG��]���	T<A�������A�3$�����*�]Q����~hcWx-e*aJ�cB.|�.X�F$I�4��]wÊ�xT>5��Y�gMBI~�)����� ��~{	��@�ywz�c�h���:�<a Va�x���������h�M�����+���z]J��O0{��h	�����M>��S� �0���M���X�X�X�u~�C���7^�v�D�-J8������@���)'l��é�w�It1��BmM�8	� ��Q������ZNL|U�U0IEih�Kv6�v��dR��o�{N����ƃk���^��6Sݙd5yD ��v£6O\
�k�M�b�E���.��=�T�R���γ�vD�X ���ɻ��U:T9�ft���h����X��*)�ν��߈�7���}�W�1�>~]{
B�^!,.B��_�*��j�#Ⱥ��ft�2*�����98�M��+�n���uM1J���5�����h��B}�ԍ%5���E�����m-����d/��&�4���*|!�����}�xv���d�R䅮|d��=�
wj�:Č�uQ/�V��1�L�p�� b0o�����G�ݝ������S�q�����YOj����Z��O~�f��|�s����&���;R�^�\*���q.5sZ�~՞''�B���j�6 �quvV�?(0P�s�3�^����]������+>[�j}BZ�3aT���u4-�޷���}�=�X��@>�y�+b_�W�=�[W��L�l����� �r���t=nW�ǐ��_
���͋�F\�aS��u�����̹-���;�G�8K�5e]�N'��
�[��fe�ZJ�6�{ � ���HW���~�}S�G�a��]�v��@͑�����}5�d���,\�/`��A��g��Zn�4yz2�q���Z���T��_�s�ш� ��8���Vb���䕡t��p�̹0�T��f��XU��O羘����<>�:{j"=7��r��ۢU����&A�N��_�Ľ�m����#ǃSlO��=��6�-�/��������g<hl/����ݱ��4���YVh�b)g)�������6�����20qd:�.��Z�J�*qU��o�,Zw�Se;�&�Xn�d*�zL5Uֽ8%+-�q����}��I�κ£4
q�J�8��6��3���f�5-}�{�}ݜ�f_��� :�ϜÐ��"M̍� �<����4�(��?�7��<�o���N�O�(Ȥ^��;2�	+:��c��i�[�=g���*$4g� Rq�M��n;���gu���u�1tK���1H��,+��#�b������nzp�n��Wi��q@	�g����V�������.��/�Xh����[{�H��g����r̭����$0�_���������ub�C)�G�ݟ�^�I���y�\�Ǝ�Pc(<N�Τ�����=Q��`�(���@9�^���}>�K!_�^�PQ��m���k"����ꯃ�*��D��c���\��}�zQ���Sc+�@ �X
�_�1��qk��6���u�oyU��k�tN���~�)��Ѵ��/l��Jʛ�L�D38�,��Zq�r�lE�i���ʱ���\����v�S �,ED����>��sz��°���������>�@�� @��k6�}��2��o!�\�yO��3�Fr6��݇��~ͧi9����_�5�Ɠk=���}���L$��i�Xa�|ݟ:�:��Y�����wֈS��K�1�KBᘓ��.��,��D�D�J��}l�g��'q:�B�Q�	[��� �����y��x:�o��K�5^ۭ�N�h�}1��΍���TQ�歙W\?��s�H���Կ��_p�q[�r#Q܍F���$�u�a�������;�N�f3r�"Ԣ�3����dn��aY�d�3�df��¾�s���Q�e�$��	<��x\�������P�n�N;v6Rfsn<�׾w$/�/]~ xb?	����������8�m�$��������b�N��"uY�vy�3;���� ��Z���G��$�OԦ�AM���(��8�y��e0��槷[dp��w������t������F= ���K�׿��H�o�)k�#o��I��z�}���������O���ei���!���*���ǁ�
� 	�"+�S�)[�Du�=��g6֨U�w[ �S BկR��i�
�����gC4�d���O�p��4�����H�x@�u�o�Q�����p��!��R�t]�L�c�dňG�QP �hL�� �فj��K�z�X�/��|m��3&қ ��qs]櫷o�#<���l����辢{�j18F���	����u��R��M�6Л� ��)K5���˽�q�U<'�ug�;�@K"�\��Q"D�8�~o�kzHH����7S�r���^ �&"�#�c'�H�Ks`�
g��ч�.7ن�.��c����4fP�c�"��GY���b�gU�����ݶ�aI��Ĩ�~ˠp���G�g�1�(�²<Phf�ǹ:>�X�u����H�^�t&���(Y5o� �����}�Sޛ+���7����`iZ�4r�*��}���Ɩ���@!���٧RdhB�BU|��i�#4�m?�ιѤ�4�5fue9��fnK��
�!1������܊��K�>6����X:�ހ�є��vF��q���N��;���(�3r�f>�e��#Efݣ�t
1G�8�6c�%{T(��Jv`i��7�,��39{<흯#}�(��Am�1@�Mz�%]��G3]\*3~����./!��B�>z�֐�% Wg���h����1)�w0N
�Q���n�>����~cE��@�K�|����S ��/�R5�A'T���J.̤������Y'f@��f2eBUy]ӤL��nE�b,�ދR�A<kt�:�WǨ���9���� lU9~���.�Lu�S����	j|G����}��[`죌ټ�QJ�߶N������OZ�1�r��i� ��4�Lplc��Ԍ���6q�'J�ò�	Ks�پj�+˪���=9~k�?�l���J\Oݧ�-���r��f�,�HW8hV�:�R?�����@�� �	�
��T��Q���ؙ0ft�]�~P�F�:Έ�l����  j�B&Ƭn��r��۵|��D���<�6e�4�H�k~�F������H���A��Cv�bx��k=��12���������;�7�p��<�*�Rr�\��ΩNX,�E"A�]�Ӊm�C�Ŵ\�x}ʭ�x�Ֆ/	}-{�noYY�5�����*�l�<c�6gQE�Иy���jTt:g�8~�6^����4���Q:=2\FX���S���$=���]��d��'J�= �,
Fc�}2v_t	쵩�U�Ll��v:H����_pK.([�r�#�0꼔}��Q=�n�=߾u��4T��s5��U~v����dR����/Y�Q��#�ֲ��o;���+��*�>y����	=~��eB^�&��B+��	d��C�W��ǝ��ϒ��!�탼.�����d���S0����w̨[��� �v������ܒ�Q�B�cwȫ���ޤ�֊�#4c��(�FH���el���uG��5[���I��֒D���q�T����Y��z���@�[�G��-�ט��_������=zD �5��*�u�=��8Eǉ��p���M��Db�ۉ������I�)�Le����y�E�64�=8�yJ(��[���۷��IIɤ��C���MV-���������HU�.-�ح&�?�9'8���!�aƎ��eң�yY%��E^��ު.鱾�;;Y���+��q���ٛ0��".�x<a�,�C >��%{�M�?|e��Gɂ�aSܺ���k��<���n��� 7ng跄�G��2������>88oQ�cr�Ҡ&U�p����T�
�.��W�v\�E�T��=wR���ڴ��Zg�)���Wnc��/��<
X��Sc�g���p�[��0�y����T����ը$�K�ߖ�,��?��^ܿ,J߫*�w\6g+�}I
(��@+E�覍��Sd?����r�K
>s�6QN?���q7��Y�5��k)K����T�9?_��>Aq*���^R��˵�CL}�Rm4���@o"y�7� #.K��P��+|~1hŹc�+���&w%���u/�&�� U��8>G)W�����Y�1��_�s%P��˂*q;_{Y�f2E�K�Π��Rw�7+���~Tz����� 嘝����h%S�3s��\�����oS��ũ3h C�;}�a>�_���a,P���íBi���������+�m&B��K�o��.��[�k�8�����4C����ɚ�kL��O4n0�Isݜ0�8nƓ�C[A���A����Ez�g��~|�Z�����}�.@��������G��ƫ(��ᶖ�$x��a���L*��ӿ)(z}d��Pf�����[�y���X{��0� ���:8Q�	��Ѝ��Qc�oY����g�t�r����1U�ַ���f��<8p����� ��8�}v2�|�����]jj�Ǒ���~�O)��<��N�L@��ͮ��מ���`и�����X]��\T���;�?�b���l9� �XB\n�}	�ʇ_����ms���9���J�w�s�7�sss�UTF��U�6�w���Wmw%�ɮ�5��h�I?�c�]в��ge�N�s{��+���{�S��2למSQq,�f��¢�]kkv	#���'}:+�^5��ng}B�Z���cn�8������Y�f�]=�HJ3�Si�	}&��U�&����|�;�܏�n$R������Q���u�������j��	4!���ZKbJ,h�3�6dh��ԯ#�Q�Jk�Tws��S��
�hc�Zq�x�m���=��~���G>�n�L��G�z�y����6Ǿ�s��):���:�����7%E��p���ߙ�ߊ�¥��B	�G���9d��c��Db����;9UJ�7�����3M�y�Jr�N���h�\����-ދˣ��*3����ѝr3����{��C%`�upS���1��)J7��~xe7�X���Gu�����9�D
�ۻdڞ9$������T�H��`b���$����o��������`����>7�15�P�{y@��W�Oxt���� �S��g�����_�)7�����I�{�8��(��";;a��Y�A��ߗ{��q<eJ�/o8=iu7��T���������v������c�7�οMe�qsu[R9MG2d�yB! ��M5�#������v_ �- ����1'��=L��y���[@2���ꍪ��OW(��n�X�8�F��?Jc�of�/2F*cʜ#�+�T���K��M�\��>�|��;����CFK�s�����r��2Պ���~�>'p�E����!Y���ڑJ�W�a��ap*uI��?GС���0��:�8ݲ����љ�c]�8�s@�?��b����P?b rz+���x���B��T�i�~
V�+��m`�x��~�KX�|��DY)�^K�'�tQ�/Ũ��h�����;���T�t(n�A�����c��|��ԫ�x��'���n��+�b�8nM��)����G�<�ỵN������td|9�ΝQ�Lх�29zC���궎�Og��>�>���q<�7���g8��O5	�qY���}������{�)�k<����"s� ������{#�Y�-�`\6���u1=���J����9 E�F�&�d2�_����k�ky	�����b���pt�8��pc�����У��A4�����1U��O�"a��l�����"��Ν��Q ��U{�	q�9�b)�;�����O@��=�.$I�c��,�	�!���0�~%2�J�j�>%��GL�_.֋��G�)�+�hia���s��+$5�ɵ;Z��(���񪮮��ꞈ팃�M�mN��*q��a�K[����8���&B���m�G<l]�33y���z�)ᘚ�$@
���[�ǟ>}z�
#�jp��B�eX���9k�Df��;����"��z��Z1�Y�gf� ���	R����*?�����+����]��P|8� �0)�`[��/vz$�jK�띍�S��궷�$��T�A���J�w2R*�ܭ�-�8�T&P"�
��v:3�4v���契k�w%���*Rv$���b>����U;e|�6������MDmѺf��S痼]W���?����|���;��Q��F����&���b.�}Hr��e+���(+���H-6�y�������jt)�a�1�I�x��Nr����y��r�2�
�l�혉B4j	ӧ�A_9�%}M�8"����b��S�#T���� ,���0B7S��R�K�x���ԥS�m8���/�2�E~���������B5h��oa����\a����`'������:�^{x���@�����f�����L���$�*-�V��'��q^:�y��ϵȠ�E�Κ�!�����6bQ�-%�Z15��aY�ʝ�E�������G��H^�ɫu���u�x����K77 ��U����'�%ee�D�H��ӌc�i��X(e�?$m:z��~�6�g���]�cH"�W"kM6;:N<m�<1�	9�\E!˲���w攵�l��>��|L�&����������sǯqc�3�U���@yU�M���R��t 7�Sn�+Ԥ�J�A_�� �v���`�p��G�	�潽��)��w��IdGk ޿�tgBo��B�$�I}Rl�
��K��$=4�2h���)�u�����][ ���w�\?%eK^#�=�f����댔*�}���\(�v�w��Zdl����O���U�/8�խ6����=�2�&�l]X�����W)%����4K� �Hw*Kw�
+]���*,��tJ���H7�,^���}����3'���߈�zxn	������RC��%c��c��p1�å�Pfط�2�Z��nlB���kT7M&�XY�GFN�J��_a�����k����Ԟ^�r�R6U�{<�&lL6Q����$EqI�#G�Fjv&4�5" �R�ֺ� ��!.���J�\X�������fN\���:R�(��C��L2��r#�tc���,466��~�}o�4޸�ox��sXo���P�3`$� O��<���]y���&�A�!H����[_A������8���x�Z�� #K]',���e'����o�kZC��ZJ�٘�w8����f��®��f�fYM�S���K���7����yծvF�C2J3����E%>��Wc+Y��h��>�Va��耡&���7�����b�R�1ӱ+ �R�>s�pP&���Pr�DX�h�<q�y0x��LNrW��v_CV	�_M�^*)(��bk{&����V|$����:�{K����:��屄��7�uҔ8^Cϭ碓�	�b��[)`|!A���g}�����^�F�����^��w�v�H�sK�+��z��ǭ��@;�D��|YWW���Ij���T�����	�[���sc����V�����;�׾ڵ����=��Έ�x.=��3P��O���WG<����?ZY��E�S�!��؏�O�!]O^nQ�:��D��^Y]]=L��T���_�܆���L�0���F��٢���(�L
m���K��>5�j�b�i��(UV�$m�k�����Z8Ԕ5�#+��l�.Nqv���DU�bSn���a�%�����`:v�����5;	�����(�6����'�}�nY��;��컩N����~I�~�T��4i-������ȉ
��W������	�S������>�4~>��:�g��:��˵i�29�"έ�R\4�#��dش�D����)��S��V��fO9�L����}�3r7�2w��Ja����yY�`z�\l�����m��4	AS���Ttj:+=|�M�R̡2���k���ķ׶�X���LoG�Ȉ^`��T	���Z�o������]�ñ���ӞG]����W  ����_Ѥ��W��^�J?����*���7NS�[%�]�\��D��;5;V#
bꪜ�~�(�S���R��~%�(�t��V��[�L����co@[k�J[��Qcf��3�s��R���=^��ՐW/^��/ԇ�įL�:���9[��X��-z�T`��Q��4�F�B��/
u�
�D̳@?C˜� �ٻ�D�$�E�r��(��R'�r^����sE ڪ��G*Q��۷�#
a�2�)��Z�����(^`��鿴�
���Tttt�s	e��å��W��i�IFbA��m��������N��獆�=�fg�:y��T�����hh����s�]翥���=ޮ����7���.����}d����y����r���z˗���K>	�~ީN{ppP`�:g�z�@�oB_9[j5x%U��	��J'˟�X?_���e�:2VN�}����ff����^��W������#�W �1G�����r�:a��b��#p˽Mlp��o�;�}�r=�#(H	B$i������
�ߺ�;�������e`
�?��L2Ͼ�!�/�:t������V�4NNN��&���R�A��\��$�PL�x��Tc�����`�>O��7_N�GU�*(�323�����\����_����_��5�oJ]CCԹ��]##�`�����W���S�f�o���)o�h��-��H]"�+��KH�?�u޵�������O�����]cc����]==��^����NLL�/�W��X��t��EhtDDD���u[�薌����2����+qqq�[[Ҁ�⿅0Qd*{l.����GI����}�
hxf5Rnׂ��u���f�ꎾ���֦��`]}}��/�r	(IeeB�Ô�l����􎯒����ߔ�x +ۚR����{���߂
o�����7˱B6A}}}fffQ!{�Ći�X��Z�چ?&�
$�q��&;��Y�ntt���b�W�`2�6775*������%����gZ4���F+vww�ݑo�� �vS�xp���qR�S�����-3��3������&��g�A �B����M��/t���|]�i5�qN�}8������H�� lH�Gh�ߛ7�������#X�9:�oni����(�Q8�6�=�㷌�o �P�o��Fi~�h��_�ffi�.9bт�z���m�V���Xn��� 8oB_�Gh����Է�����jr�r/��74J����-����cNɩE�G�n��ۛ��$\^�[C�O�Tݗ ���p�wy�4L�1��S�t���IX�^���.����{�/[�6ek$������rh��$m��?.��Hȸ�fB<c�"j=: )��AIii�S?:J��կcZ�x�	e&#���áW-�C�����〹�ir5�<�$$�ہ������
3��k�!�o�8�̓BϝU���C��-��<k � Ov��vyɃ��X��H�4P,�}�?�����7xs���������ۧc�������������i���x���%bb�u��%E�H��J'E�[��h^룗�:chsʯ�T*Ǌ̗���b��D�z��R�XT&D��@8`�L����-###��Q� �%z����}�����	��;uA �Kz��g%�*Qdgw&����!@��1����OEE|@a���9�؞O�q �,�۔z(�\�/�*��l.�I�U�m�ID/yt;�*��}٘*���ݧ��D7��od��y���N��G���������ʆ����o�F��w�H�j8dbBmLf7<�v�8��j�t�[B�5ZZu�H˽9������P�I�?�.�y� ��0*̀'chH};��p�HrW�f��`����v��V&��az�w[_u���<l�������ͧ6����\\�J%}�C1�����?��l��*�un-:���1
?�x���

�4C�hK��x�.��<,�uI#�k��b�A������.=�zooo������GW� ���l����U:e?+���;�+�Y������ �L�%��n}'1�����oݒ���ѿ�h��S�$�PE�R�֎E�Π�x+6dzkOUI���C*}���㑮�UXXXn+6h"�RaZ�	)W��9���4=ʮظ�2����B��CqBO�(���x��{���->����"���%%��F������ �+
]�	��Y\��x��h�_���n�=�� ��d��*-��o��H@�W�$��͸�쌌&����z������]r?9T���{�T%L�l�CP�0��\��kk9;�g�?�)��}�S�Y�!ƚi�W'f���x3N��6�J�ffgˊ���-�6�8˰�'�x��4��x�}LM�.�~^��CD�TVV�H�7���^߻{���K7~��L��xv���R�Vjʮ���5�I~ܧ@��a]ʿN<�ƞ���N�M6�U^��j�E��z����x1-�mKK*���[��G��	�'5�G_[JW=co�g�קv���6<k�m<<��=<t��$�\�ӹ~7���CU�x���D�8���1P�D����͇���><s�Lޒ|Ł�&}��#���n�e�S���@���R�VS�Q�L9l�P���b����~�k������F�C�v�I]���������z�[�Te��˩����� �9ؠ���z���d��0X.SfQ��Ж3�4@��LW�(0��p�4@�n�Ȍ�	���w�g�d�Cz���!��.R6MM<թ����OQ1X�m9�K�D?�Gn�����dQ�搛�;ۋ�<�뛛�����e�X���� ������vv��\e���@TLll�#&�3u_����H-�?����~���x(s��H�u�J_�OC��|��������d�*h\,lJ8/��w��g�a�w���V��nu'q5�g��d�����b����� 7������֞�(a]6���]]�7�3&/󱜾�F⧹d���-����b�歆� ��Z�>>1���0&�$���
|zck�ʝD���W�V��.ՙ��3AH��OE�-))	I��x�ߑ��.�V����Yck>�600��^�u8����5y)�?��	�����"���]A�������������𤨇��z�]>�c�27WNc��=wj���Q��>NU�ߖ��m���L�C�����8w��͎���lK��䓳<j1�Y�㣦�r�AMC���X���amY�eTTD� ���g���1bf�.���8	�������y	�O��z��d:Q�R�5�Г��E~z��7h��M6�@@� �V ����|��n�ؗ���sf>=���Y�^C&�C�%��W��*7d؉��K�ى^������S�[R�XpD+��?�K����<M��9����@�Y�)�L����������Mv��F�G`�c���:�z'c�s�tR�i��ữc���w�"T�Y��Y+5�vq|$�uư��}䜋�@W����{�������:��#����BBB�yyO�g����9���g ��2�I�S:�P��ǹ�睊�c���Ǟ�ǯ!^��_���V�Xՠ�Tˬ-~�!�yyT�U.��¿X1��H]S�j�r�y�W=��B4(yyٚ���r�ڍ��-���ytؓ�P� vl��4��c?�
|�D+?����(�d�LI�Ǜ�E�/V?�R��!��=�����}��h�8>��tP%|�x;��7�"��7AЅ���/�T���.�8I: ��E��$OB,��ؙ�lZi���1��k����F��Wx5,HHcz����jd���f	�����Up�0�w�n� 8���dE��2

���쇚��BDEá́�O3�u�.��ﮜ������F��tp�p�X����f&��|4�%�ij
��0fw�x4�]h��8���/A!d���~� �DMQ�r�Y����`����i+%v����u��d�q	љ���s�f��-:���:�[�?̥�@jME����"�b�е���w�#.{r����?��J>>�.I���P�q~��������yw�?����5!&;���^5\z��X
t��G�J �?\u899�99U�o���߷taqQ�����.���I�1�����;�p+�T�M��օkྼ׌�������d__�5:��� ����@)�@)U-�,��@����Ja��YUUî�I'q
���F�Y��߸;+uP�G�)����M1��/N��˷�.4��Ns�w���@�'�=e���=��٣�{��V�<C�k�c;��؎j(K�04a7![@�R ��Y�	�J-�'��S���A��_����ZX^Vc�Mg��c{���*9��aq��j�@,m�M+�����1q����hp��n�^�� Hmm����rsU��31���0�ZXl�j���E����ϯ-���d�b��ъ���[�ŝ�,N!������R��C6�.  O
ZZkFC(�5x�Ull ��b��^�g I���C�b<�v��ٔ!�2ꦎ��"i !���I�� �4 �Aa�?Tb�;:�k%h	�b��Jl�3V�?�v�3>���e�q����.شւ$�m����D����!# ���1g+��7Sɢ� �d>��Θ��ɫ�3I$��c�T5�RE�u���	5���x ��[M��uT�m2�� ���R�x��V�(e��ڌ�<TUWϮ��JThr�hS4����xg����|���I�~�r��P�MB�����Z���+�v�R���� ʚo�Y�^qԲAU�iƚ�}���q#�C6c�XQ�舾'l5����� ���t��̥O���n��@t:�	����OJ�̴4)�����W���j���k�dl�����-��s�v��EH#%��
��Е�)a-�`���X6�i�-�u��z���kHb$�PH�hm��5kcl�����Z7zp��<R~8:�����H���)�^$��`����:����*qZT���q�23�1QO+�s���9��I0}<�X�[�x5��*swn��mw��j�W藉9 7`��^������%�^�n��G�~�9/�h��|"��<�*���N�%Tf�A��.�ӷ�N���G�EC?^h6)Z���B�~������x�N.��եH|钙��0KZ	�ĵ�N\��#倇�O4�jw���z�0wuIۢ��m������	wK3��d��� ��r�s��j�U�&'i��VB��=}����y����q��=������a�v��ʘ�(>|���lUs��| �����ѭ��B^UUՓ�n�R<ğŧ�)���a�f@�ݜϢ 7�>{�yT��f�w"��}6�g?�r��A��+~��C���L���~�:�
+���;7w��J>�UyR8�YA� ��Ԡ�ߌl� =\zm�S��r�N������~Ȥ��6}I^z4�֡���U�*��h�!d�r3q|>�t�K~/�Cl���1c(�塿������@�[~^�ey?WFwUdDD@n ��N�MM8V�O���++�zaCG�^^5��H��?�(�}�Ձd�v��+l�Gf���:���u�i1^��g ��6�Nɤ��Z��B�D�خ��5Ͻ��ƫٴ���FYY�B��Ѣ� q���b�ٽ�Q]�s��M��ސQ���B����g��(l��2��:N.C�^=N�c/P��Y��Q�BN�{U�q�PìA,���q�2}�@��HT
B_KT=�D~��?�����;p�i؄p4�=��D�� A�Id�{�����z����A��J�J�c�5Em�V��H����פ���Y�B���Th!=w���ڽ��CV��,zw�_Q�����J��ڠ|������KY�Ŏs_�<M�7%�\��k�`�����Δahxr�(��?�8��r�?�`���W�S]H:����t��()Q��a�G��Q[����U�\Ba��ҹ=[����w��a޾�[4.��|� (���:
= �~�;V$/ۻ�]���Jw��Lށ��jjF���(�ԅ?�vE�� �Y��G�`vYp��(.�wk�M	��;����P����mL��o7�E%���6X
�(M-qXm��?rwj�๪"L��F	�^�9��C)��+�V��ҁ������ggg�J����E�~!~c���.QkO�\���}ZՈ��Z��\hh�V�2�}��~�P��M�W]�pK@�ٚؖmXb����@)�ԹN�ӧ@;�����}v�7��b"�����iI�#��Q;Z�e)<�8�Q۟zn\��/:���gk���6y�l�֋�$9��TB�-�U���.cOY�m	�O��j�IUE����^�.�_g��:;��3�k��7�j�Xk�I����P�#����Є�3-	�W�?�G��s����e�U�_�!z�\�RT��;��GS/	;}p���4�N��q1�YUg�r�����������wc;�fz��\��*������m5��q�l��������	���9� �K/�	=[-�m�RҾ�Ψ��B��U��W}��E$zGΝ�\,gV�Y�y����&��t��&����� �V'�	ș����v=����b�ϋ0T���Q�;�Ui}+��YݵCqRg�K
��&	�Y�^�9�]�s�Ǆv����H&��`�"w�kV)f�� ԅ5�j����,W��WP��Wt	���N=����˷�m���b�g�+��f�|�t���r��(��aƸ�O��v��ѝj�;81|�
gB}������ùSV#�-vL�AW�ծ���f�,Uj��`�%����7�A�r��JE6�N�P�LEk�𪟡f�T��L��,A�d��5¥p���z��^�2DnիM!�2O�%J�=8˙͛��H+㎗����[�1
���;��5����R><1��}G0����(�/	�+AT���>=�����s�B�����lf���fw/n:�\#9���-m���PZ�9���¹��%e�qf=�J w����C_v�S�;��k��
�i2�Y&K9wfګ��o�Չ?��E8�n��?θ����ֿ<�M�ƙ'��A
s�Ke����9�գ�ͰF>�<W0a���n�����5ˍD����!�=�7��}4x��Â�]77^�.��ݚ,5-��z�Ie��}:"���)�,S�A��biQ�T���oD��˹�b܋gp\i�6��}���&�U���X%�٫����L���B|]��fK��R���Ɖo)�1jѲw��<��\�s��w����o���v+f�1J�e��!3���[���b�A#gv��D	��(�� g�2�$/~�r,��U����e�sAS���QA��STXԧ�\_���I�^�bկD��K�F���K�W�?�
b����k�y3���j�z�~\�A���>1��ה���vl��ӭP�U`�B�2s�8��GLӶd�<7���S������L<�.�P�9`4��P��wd"(" ���!��2�Bh��~�����i�ͩ��Su�Aa�2�7FB:�| I���̰������"�l"Wl����]��9�:���rڄ�r�Y��J�ƙ!!��g��z~/D}}'70oC�)*e�;*eK���|x����O`���w����s:.f�K��+�ul�p�i�c��zu�6�}��O�td#h����+|ٗ~X%��d+9��mG�����T��B�J�� H��]��/�b�X�]���`�v�=�,���t	ۈ�LM��rC�i�}oʟU��d+�hs<{�Ԙ���R�mP��aZ�v�\�����j�z�Lq�!�	@���T£�fn!۸1��G���zr� }��_���s�rV�>5%!��ک����w�{{f��W��H(s�w��$����E��p��'��d"8rY��S{�����\G)��{�PKE;%�1���.*�<��!�����/)<�A>��!�ckd-�+�슱������m���*--?�N7P`ZXY�ӝ!+.5L~C&V�;%��:*�Uqf�a� W	V�fiQ�@��jB��U���H:2�����Γ5��1�V;W��*����	�;��p+��/_�����;G�#&�·���#z2�o�{���&��ϡ9T��¢ڣdE��*�v���KUّa�#Di�KRj7h),�5b���N��j�o��e3Rj�<ZM�\��勫��#��Yw9麳�.]��0��~��:�����!b�z�"l��"0g��Kɔ5�9̻��,w0dw�c���3V��߿�L�^�b�0Z8�	=�yJWW7�������N�Q���så�s=�gL~g�Ɍξ��t�����D}����kS�w76@�*en�%`�	x�3��GX�:i�AӾw��Ҝ��4��f����ہAA1 o�Qv=��0���{����l�=�F��55�����!q�g_10��-MwS����"?*��B(�i_�g��?�RS���yS�u��Nh+�۵��S}cX]ɠ6�i�#�(sr�P��tHt�/o�3Vā�4i��U�Wk��r�W`����T����g��z\�&��� C��UQLG�Uo
8�TK4�I��aٸ��b�����C�|�2ā�C�{s�@N�=��P�;�k5z/Nu4�-�?Si���W�C�f�r�"ʝH�z%�?[F��;ܖ9�d�U����  �}�|U�ec4�;}s��NҜRj3n9����x�A�I^�v�kI߫gyb|�BG�yI��if�ߍ�)ֿ
�E��teRl�����s���f��
�ْJ�S1*]:��{.Tk�O��E�ͱ�]��Ra��M�X��v0����zd#�-�������R����밴�_6�P�^�����InN���6�����k_��N%~�d�2�HN�MʦH��MW��M��.c�\�(	�2�;��9�-?�4��7?��a=�(*R�#����\��aܓ� �o��9����m�[☠_��=<���D��)��z8��p��~���Cyi]Na��$��MLM��⭤W���}C�mq�����MrC߆�\Ŭ!O��k���	��#�Сr;Fy(�W;ڒ�Ld�(�PP��{�e�	)��Iȉ�~ۏ���@E���[��TfH�������2:NOXƄs�}�8s�w���l�H�C}��9,u�����yi�)伂-�(�	��z|� ���*���e�t0����d�����5���4p>_;����c�U~�P�)N�떋[��q��*�m�v0������ϋ	���p/���2kk5~j�t���ͬ�"��O �JJT�+Ia/>����MI�WN����˵@Ft~i��q�Q'o�OM����8�u���p�SւA���ͱ���?.(��;�3���l�����U��Q��t.������<�+�ic�ذ��VVPNNN����n"����7��|mn�����[��Ťʝ �ாL SM.�oƩi"�����P�)��x�8����gપ)m��;�H�*9���ҍ�v��3�����0�%Ҩ�<=��W��Н�;z�t��c�r�D ���v����+��-���[}�
�P��Pf_4����|	���ܷ"]!�ޕ��@��\����%��<s�,�܎�fFb�J��2�cu|�� u�\�vY��9~� ��򟾜�Q�[U
��V��Y���c�,�q[��ݜ�vl��I�1�:��y�Ң�U՗S��z�b��W�|K��v �>!�)h9�l:Bb����Z�U���|,�p?�'�_��Mp`#)d̸��Gz�4XUR +�wC]`2%�������"A��+�eJ�x�;9:��?��Va�r���,��B^*�����"�;?*,ꉱ�v$�ѭ�7�M�h�D��bh��L�޵s�zSh�2y�~�ah�CK:K�n#)�~3nͭxǋ��>?o�;��(g��u9gx���-���	y��j��$�iiR�{i��FJgΜ���B����Უ��ot��>|������Y�I��#��GLL<�1`���dIKro������Zsq�����1&��͟���IM�AV�ep9���oN=�F&8�V��K�̖��v5�v��yl�Q���%xOgk)��3-��,�Xٱ]6�gZ,���Ιm�]�W+���.�)���?��UURJJJ���b釫Nrr25H$Q�G��S�Դ�=߿:�ܷ��EEK+��g9��nL���� ���b	1�[;�D���aUar�7�����-ReIW��-I����Y[�|�p�s�sA�E���R�-�Ĭ�F�8I|�S�G������x�>N�pd=�|�&!�$f��M�]���V9�r��k��!c�[�Nk�l����Wr����S�uvz�}�+�*��w�Pl{�-6U��f���+�	�T�Skk%666dB����'��W0]1�����RH6V��P�5q\I��z���|�F�\�����_��I��>R�X�"��Dr,�`�/B�����Zq&���F��`�˵+��i���ؐ���I���/���NS��-?�GgCϣ�7�K�e�������8�z%�9O.�,�а��C��@��4W��5Q}�7�rk� #�@;�y��_�A��+!oYx�j������gg/�7�s��ue�	LF?���vL�誫ke�!W���F�K*l�d1�_<\|ҭE���y����A�{�����H^��@��'li�S�{�t� M�F�{���+�/T&6 ���:V@0�/1���IݬdO��k���� �'�'�/�^-%�q�s?�����J�=�����xWT���g]����YV�������a��6�����A�b������#M�Z_	�c4�!X�.�U�)�M���)�%#=g��y�ˠ?Z8qȪ�o�l���0|즗��.��J=k��{�7����~n�Qr�5)sɹ��g�U~����0�VlN8��m�X�Vb~m1���謸��0���r��~N_��tj��&а5?��{�)���*����%^�&y���	�ڤ�z�WJV��%�s�����o\X�ٻ(�
$:��Nhfrˊ���vB��w��I�VU�zx햍��nH�5��+C�շU��Uc�����Z�]��$��<\&\"Y�h���Q���9�2�󬮎9R�aRI�=x
��c�]�-"_�q1G���ʻԮ�O=��)��#�	R�)�*�-mU�1c����07k�T���⥒$�o�M$��պ�)?3b>�?U�c)���W+{T��L L�?��}�Arşrr����,�����6S�{kHG�u�����<���7QT��	�r��(t�x@c�.��6mQb�������Cc{'[mB�A�pHs�J�G����ZӝpF̹��U"b8��b�I�x��s�T]��0�|u�<n.z~�+ɂ�H�
[��c�����t�
-^ڷ��I=���RW��/	��3��h�n_u}ǁ@}a��a��1_S�{�%V	�>�^KꤿV�x7$�KM��]#���#S˄j�üeHs�s�˪�� �&+�B��N��d�;��)�Ls�Z�ݺ������g}�����&ӻ�ɠ�d[�Ļ8hO^�h�]	Z����!�Q�4�� ,7��s��h��P]kԷ�10����I��y`j#��9�r`�,��t�7��u��Pތ�ҺV�����#�@-b&!~���йoY>���t�U��vp����\��G�jv)�Z[a��z��DI��=����hT٧!V�k5}������o���>�3]�[d�R���qǢ����H��!�c�քKb��t]K�V�:��`������X�U�1���T� ������"�+�=#��ڌl��䳧<a��Y�^����A�-����ړ�E�a�}�Ӛ�����%u����ݚ���Wo�#wEyN�[�a��7��]�l!%�<���b��TZb�#���o�.y�E�+�.~��D�Sd�d��O'vY1W���_mIa���	��T%8�U+#��'.#�F��2D�U_A >�4�9	������rh�\����2vZ{o�4�I�U��G0�p ���RHʄ+4�VFi�A��ha͵�s;idFZ��1��Z�e�v�q���1?}��x+�!����}����~JUo� ;'B��~H�?XH��x��pJ�=D�!䍢�h�h0Ԛ��ƶɹx��!+�ƚ�%wtS%p�u��ϿU+!�J|��튍���������������tMa���KZ���}40�=j�����%9h*�x[:c��A��d/G1=/�RZu��YBݞ�,`P��s����� .���98�^=KP��H7�C�_T�

	����Y9��7��Q��<ߗ>>H�ֻ}�ұ�ʹ����A=���2A���>��e�:�xt��Ѕ�8M���D���b-�����ț#�M�&&ٗw�ᔼ��5��,��H���}�I������s[�f�e��Q�|�*��;�6�;6���	Y�ܒn�D��;�
+�
��х��.V�}v���0w�>�Z���RN����p��2o}��+��ǯ���$Ӓǧ8x�e�-42^�-��N�9�V)�����s>^5ǆvk"�yz�k�]xoq1q�1���O�n�>��g�J������Du���$$WD�E�5&7<��5�����Q�����V�.�s�й��h���h���~�T�흣�j�ru�e��;�������ZD� �a��Gs��NG�鿖?l{;�$Q����#Ӓ:T;덾��Q��-��LQ�����c����	+���LI�a9V؂��+�;���>�C�vc�Z����~4d�8)N������������=��)�d�8���0jC�M�?^��+�ן��f�U���.��"%�I��QoYi���go�
:7H��뾻
I�����Zl�� �oJx׺����K��X��rg�UU_�Ғ�>���@(�?B�2��k:��B$?G�\�6�+���ь�>�N�P�c��ƃ�;Gpޠ#�ʵ��B��T-��>Ii%�����^�"I���=]u\�Ú�ƞK��,^cq������6�v%3H�2�i݇nZ��!��DK���]j���^A��ъ&����(���CV�����e��U���E*˻<V��[��}����]n[:%-����>n��E����$�&!���8�x>>1~���:���ײ�צּ|v�m�;�F�s�G!Y�A��o�m�gnX�h		n~�XJ�@:���n#���,�����~��ò�W��:~ó�ٔ�~'������g���Q��>9�/GӦN���ZWn&|��F�\��|�Ԃ�sT�T�2����KI����������K���B��
K���:�wf������;]�d�8Uai��(ϸ2+�w�nϻ��/�fCM�e���W[f�8w�fZ4�l1K#&t�S�v����2�^�59�
�0����ܱ�Te%1A'�T��e��8�M)���p�f��i訚ʪ��3f��n&��͘oy�!G�����g����T󦝇�myD"���"7��:ڻ��q¸�A[�0��dd��
���P��e;�Z�*��T�pC�f̓y}���A�M,`�D*��s��!=�%�A�<��c�O��1�Ru(�5�����'���*J�й�MB�>��3Δ�B�f�%|,i�PR_Q��9��sY�NǵG鎋�_����he��B���H���>̤zw�����+V��(��i�Ӻ��2�Ў�۽�zp�GV^�T����)��!��іS�,x�1E�j@ߚ�	�I���ß<�.X�����u�RvYx�ɤc<��۸D��QY��N㼆3���ÕlY��
�t�{p\܉���#K0��kL��
�n���17Ar�ҹ�Z.���'/77#M�����aʴ=ެɦ���_p�+���m���k�c��t˭�����=�������F���8� �t@�O1��te�
�#83|B��څJǄu$�����
j�eX��U)�s�1m�4����ؚ]�E��|p����:�U�,��X�氞j�U�K'������+ʎ���?�6�0'���	�=��1��Zm�x����8Q0��,@��AEo�癲u��@>���w�N�������7x��U�1�K�Έ��x�c��w�>g1e���r[���cȎ1�4r�t�u��$P.���Z�%����e�>!�s%������G�-���珛ch�}Q���m�
�i+�b��XX�B���a�i��l�oz;��,�_S��"�9���F�,jk�'�]0��f���n������ۨ'�+_�b6�̚����򼯠cYv�G�޼U��2�x[H�!�Axb�U͈<+�4"ĸc�n��k��0z����+�,��F�r$��	z_R��x�_�v;-a�i�3�I|MN(nn�Ĵ^7D�E��õSU!o��G��&>Ω�MN5�N��jkЛ�B�ý[���ˉ��iEK�Θ��O�r��T���嬅9V����y���HQ�C!D�o��^��W�?d�IM|����
��
�| Ʉ
f�=��$�_xG���Xƿ��$�&V�R�_L�b;�܉	�8�����	F�Ɛpb�B"��!Y�y�X��&O��}� ����8�G��u���Y�sn�Ee���	ۅ���tzmr�Q��(i�%}m�EoV��b ��yE�s ���so�������|��:����!]�4�l��'�KA	�:�n�3޹��R���h"�>��آ���u��k��,�zn�1 Ly�WF=��]#X��!�>Y 5��̓d��ˀƯLI*�T�Y/����T��a�\�q���6��hcI�x���=�X������Ԣ7� ��`���j��Obe�h)C����yQ�����������r�?�!7#*�U��_��v~�GA1�jm:��(�ꐾ�ߋ R[�Rk���pSLQy���Y�����uƋ�ܓѬ�Hp��d�8�bp�r������N��-�c�2H�g��(�]+|���&���d�H'T}T�U�۫w�����;A��_ԡw+�VUʺ�I��_�a��t�,�g�vDӪ��9ͧRF ���([��"�s-�k����;w�P:e�@L�x�B/'����o��3hn�,�IG�Kv;���H]ĶP"��ˬ�	ե�O{S&�	��3��ä]�:��	�����+ɭ������7Nl�����f������.�������2��z�1D�����ѻ��/D8�t��>�~ٞ-ɠY����B8�]�`�LxP9v0�9G�[���:��~JowO��'ٴ]jk7΁,ș��q(�~Ё��z�O��q��%�ڃ=�x�'N҉��%��$y'�k�T!(���_�V��g�)�r�.D@�GMգHk7�Y\�+w�)8��Q�/RUq!�<�i�N��Vu1�BLD�����_-$��F<ΝP�.ྑ�t�ցT}Tqޢ��L]����K�a��7��q�>!�6;*eF���7nF��=h�_z�U%���u�}�d�n``�Ҩ�<5���jB�u�j���|�E����"/MȮ�bd�(�"k�����|l�Rb{Q�����%K��p��[�G�H��n27[�����I!7�Zo��G�L�LI��B\$��l������������T�!�$���E���FXFG�#m�x8T�o[C�I�@c�\x?:y�C��Xf�M2����YN�cO��^N��3.�a=C�C�K������!���Tm��j��ô9���\��ڒi��匔>�s:���ºw��R`d��4//WL�^ʴf�_�Cz��]hD*� ���ԕ��<%��4ܿ	7���W�6���������K��}S�y�^���܋��<=�N����*o�(N��U�Ҍ�K?��x�s�|{l"4K4��u��W�א%j�p����v�`R�J�R�>=@#�j�^0cɡෙ\ωs�ߔ�
��gV&LD��zS�TG�����������t����\�f��N=�����1�$�=_)H=�Wyf&�uS
�l~�hl3s�lh�砾B�iq��H��,� ��q$
Ő���/��*�,��$[���?�Ye��z���Hܜ%z�{�5ө�i"�$ktYV�Fg��O�T��Oz�M�g߹nBF��<4�{v�z�p�"���u��>�5	��8e0��1_��n2gO�AZ,���̽{�<cI9Vi�@�?�B�b�75�ߧ[v������Aqu[ yyn�IB�wx܃;��� �K��A�C#�K�	��xc�6�����n���3?曚�*���k�g/y�>{sJ���u�%+��%��$��_��-薃���e�N[�S�<��
��W�����͓"(�^p�Kʨ�_���+�S#�Dth�'eH��R������c_]7O�-T`�ޓ�|{�ApW=gØx�M�~�ș��ϧ��Qq7�W�����0�>9�8`�П�y��qǴ6�\yG��DA9^��<��.�|�}"*|Y�y:�
���N���G`�k�-ז�:�7�����qk+�*��y����v���ߍ�d���"�{AY������8�j�o��W�i�ى<%����5�хE�À@�o,|ƍZg�ҢQ(FtkU��7�}%0�����aŌ�dwz�!���8��Z
�����q'D��A�:�Ur��IX��J�V���|Ɗ�;6 �I�{r 
V�j�!/��5�n��-�QQ��E�1�J~Qg�D�q�ҏ��ܲ��N��sƃW�� ���ǈb��X�e���r�c��(��C�u�w�O2���R�����L6�O��_yݴh� g$n=v�����U-]�>��M���}����u�- %�)x��ţ�u�� ^�L �zp�]��5ʛի��JH�]�j����@��ӖR��o W$}���>�;^5�A�ԏOa��j`!�-��]7��`4�b�F��B!�NG�{��n���@^�Q��Mf�Y�?w(A�d7s��fFšÅ������G��ͭ�|���~�ޑ}@��J��8��z*�e�R��'w�Z���⋱XJ�	�����-��wG��< )#�zzjmg*�?�{L��r����!��\}-Dj�­�w*�����]>U�0/X�`I��3���&�ua�xIa�C��o�v���<�(S5��9�?�.�t��U,;^$�΁�
�V�N��R��W����F��j�Ϥ*xQ��|)��N��?�#*��[4.2ɏB�m�Zt8�o
�<����W2�q���xIj�/�U��gK�X�,r ��JM����:K��4�F��7�q���}!M� "`SE�֗1PA`pCE���>�+m��s�#*�2~��ݲ	�|���}��3^��
8���`�p�����(|�C j6�O��c�!���Xa�+	���^�mU��q�c��l�6>�������x�Z�+����y�A���'JZ��ҭ{㌇�+��5�,��Y�֥��\��I��m�]_Fr�%��7 �a!<E�x�d>s;!�31��r�<�h�;�=Z柨
~���n�X��ٺ��*���p�;_ngp|_eZ�V���az�6ؠ�)�J����۶��+C{P��o� y0�h�� ����3#�t8�� ���͈ �]BP*Ͽ�s*E��]��xU�L`4�D�r�@�ԏ���A�l����G�K��'q�n>��]o�r�Pۡ��B	7��Wv(�s��;Om�ݏ+�8˫�%�@7p�}p� 4�����m�^�����?4�*�e���ϕ0����yp%����C���g�k�^ފ�8
�WAOĤ��u��QP���� ��  H�dJ�W!�_Bc�����k�'��c���q�+i$2�M黁f'�f����.֢��	��cݼ��qw5!F3jd/�����R�	����^�������E>a`��D���a %ۛ3�ͩ��'{]��~����fSC��Xʴ��%U�;�Z�}tل9n~n{���g�?obz;]-� �I�`�ڸ���<����8s����Ź�g�܄AY��_������!R�@j�b5���gK��
{�	Eof���a!�-�_K�Q.�r���gTUq���Y�lZj��	����UyhxޫwU�T��?�XV�#g�8<�v+��̆_�!�K�W�y'o&8t�T��?��	#�TK��q�Hg	�ɺ'B��)G���?}>42N9� ��� �3��OĀ��b���@���<�9r��t����oIsŞo���11��fW�ޞ:���\��}[�A���˟JR=,Prw���ӯ��}@�0QN����2���Ty��1vO�ط����!���H����<r�:[{�քe���2���z�eʣuS˶*H��/>+'�_bKU����X�?q�M�lH�̍-'�� z<G���Z��c��`�ʳ[�N^����r3	 ���L���Pr��Bd7���|)ױH�O*q�U��z�-?�o�y0���^K&��Mw0�� qe3]�foF�*L�|�*�b�Aըz}��̞� *O����m䝜(O'�iMƩ��Hʛݥ��%���WP2�T��jb��T��`[7�\$�b����Qw��Ѓ���V��%2�f��e��3��]T�}��W�D%���f���S��MH��M�ȆZ�&�����{�s^�cP�\ɖaV�pސ�Xh`gS�����M�]��N�ne "�D��PQ���&�O��-�B���ZN<��MB�ܲ*ß�#�v�X( ��F�e�>�|7�3��0鍽[����0 ��<��S��9P�v��ă0�/��l��w�ܽ�9��+9>��z ]�N6c�L~��W�K�FZ��xZ�|���G���=��������1&{����˔�_�1��<�w5��=�N9:�u�W�r(hc�8�T3��������Im�&�-�U��?�M� �U\A��� �cË�Mgy���8� �t����͟�#����?Ӗf��C��<��`�a��9q��z*���ê�eߏʀ3�q:$*���W`�4�{n��V?��\�e��t�(׎to�����Ɏ�_���ϖ��QEA��� �w���F7ƚA�N����}�Ӌ\���R�����q���Z�>�
���\ȣ��3,m�y��ʁ�U��6�w�����e����/��j�}`�+�q�ȷ�zi�އ@m��w� br���z$������"e���?̻������R;�#��=��ɏ����˫<�u$���AY��U'pa�`��u�}�;rb���N��x(��-��QϠ"s��d�]����Sg�	7�'���q{���	��rT�2�5%սx�Σ�Ev��[29��``PtK������ٞ���b&��*�%��Z��&��!�����`��tQ�� ��l ��m�����9<qD��g�����;�G�ؕ���̻�j�Mj����C~��u �����:����(㓧�b���p�ݬ��R�ͺ�պ:��2K��}@�)����5�&a��b�+�z{��v���	�S.s3���ܜ����}��j����syA@��=��<-�=�@��y95�;�
�ïO?Y�E�����rp��Z�t1�m�6������3>1�XQ�-QQV��%u�_�9;x�l�����
%/O����>ew[�&XgP�B���"�$hS�	5��v~ԩ74�<����Y(6{#>�	'�.���VD킳X��o:Q����0��ܙ�-#
NɆ�	ȃD��H���;��zs�@�|���o�Fg��'�Eu~��(;��?[�u-%�\./��Q������r�k�϶t���<��ݲ�d�Ո�57�<����[��5i���Vb�<`Wj��tj<���d�Ԃǫp��1 ��m@�uQ��� ���IR8X���T]�C�ÙEK��t;�g��d>ա"�����-�7ݰ�<K�c+�!��Lq����y�}���D��B�����<}�<�;�K����L,߰��G�Br��JZ�]	p�"� �t�u}�kw��+l�O�R n�ų
�u�~�a����y밠q>��a�@���=p�t�
��G�C�x'w�·w�L��<�d#3���j+�۲#�DŴ�`+�#�g5�1�����}�{T}J�)��@@Z8yO2�7�`�Ra�����=�i����U� o4�Fq��Tզ�:Yvؔ:��,��X��|G>�4s��BK���Axs%B�"�h�O��L�<�=�Y��@��ݫ��:����s�	6YK����$/bp��n�;�U��p��kA-B�B���t,�.��u¹o���w��;�(	�9��Q�6xe�L.%���~k�WK,���܋�H͊
`p���R g#�Bπ�½)Z��'A��P�Q�d�k���p_q�Hp�9dc��mD
je�52���_�?��KZē
�%�j$�1�D�!�����d����w���)����jT��������
ϼa�@���~��Y
_��*�l?�8��bV��\U�$D���o*�-�@�W3ֈ�v�ߑ4&�<c]�d�z���K�Q��YQ�e����GtN�U�&�28{6)�ƕ�O���y_�yd��S?�y�!���������^�%�7����z�(���6����o]/��[t|�@K]T�����G���)\ǥJ���(�I&���bZ,�Y����RO�_6�L��ۼ6��\���zH�	�~�]j��E��[�6w�	r�a|n<�2���4���E�9GΪ ��Z?�d�aN����]��{v,P�.��%�L^{c��� ���ԽϞ��o}f����d�d={���5�mM3k�N�0�������p��~��w_;�?S�␵��z�D��̫	��ŉ�cw�n�aVzd:�4�o��ñ�[]�t9�}9�Gw#=�������Ի"��3⃱
�C��V7ȯt�L�Oi����p�9�v��b}e�\���e��+�n�ɓ�.��p]�]�Z�}��~��P:�A.Ф�ZTsz4�D��3ġ��ps�e+x�z��x7c���3vS�q7�l��Qb�%G�U�C.��X����y�^�>#�?[Z�]��_
#"���#s�����;2����?땯����C����㍽�#VO��'ⲝ��>�Gw7�n�E���%e�de*i��A�cc��v��X�ϖg߉+cH��D�A�G��p���)O�J�6��]�#���"&V�Z�zԕ�����O�������l����]��7�
�M����d�|�a��I+��K�I��x�*���nY2�آ[9�J��2Z����{��@�sl�㧉�p�N�yN�����qU�{z=ru����8���Ԩ<"�����^��w^�Y�'f�*����9��ml�5�X�Uھ	�|�T�ž�l���`���e"�X�3��ن%��	���d��a�.�Ņf�H��)�ʥ)���$��	n��ݷj^BS�d�h:��Ъ\J�e~��3�i��q��?p�s�-ꊣ�BD�Ȧ��46�����:���H[�u�h�ǖ6���Sύ�Dʥ¤�kMfE|؍a��ϔ���"��u�� |��1h\���ii!s��7X<���;�vޤf�S�d�dy����͝<�����uŨT��\'q�3��hTIUt����5�)���z4��`r\�:i�G����v�����fD��cTp �~H�����m~*h���6&�
�����>]�����ŌG#�Y_��^D�D��[>���z��M��)��������ۛ5i*�太1��N���R�d�����?<��4�hI��7{�G���j�= $����r���K�n�(3Q�
��6�$��՟z99+l�w��~y��q�wCu���ĉ4��3�_�o�J�-�$�e�r��aÛ^,����"*��B�԰�T������'�]o�EFK͜���E���c�Þ��?;B�H'u��&�X���Mb�;��2�B<:Nȭ�:Ǧ�tέ��>��is���J��ê�Ņ�����T�sm~�J\���Me4��׵+�֭��D�N���EI1��|=m]�9U�1!F<����Vr�C�(y���]�jG�o�!?�k:��Ξ�?���p�l&<S���m[���ň-��=�K(l���İ}�7��#O~~Ĕz��>6�̽����(`�i�q5�~�>bW���fM���W��S6]ɺ�� !	�.��s���
�)�X�Y�D����,��EP��X�i:�b���H����w6HV�p*��O��M�T���5#�_^K�??J�X,����>����Ys�n�����o�i#E��.Ok;TJ��A=es�G�a�x���I��!�P%���&ɰ]��o�%{�� ���C&5���P�V>���j�c
)^�H)�N��P�0U�G?�oX(Y1,4���6ʌ�S��k?��HkMs�T-����p����C/�QNb,�a��kI��8������B��9�]q����HB"b�K���$y���kkvVrbC�%�[�����6�ȑN1<�i !L��`J�"s|��,YI2�T�FK;K�k�<I�ї�q
��̄��r7�{������%�����<��mc*7c�i�l�i=P:.2����l�fě��1��Ǡk���}�6O\�L�D�O8<�Κ�U/-��zy��P�|��mNC�|�
[��,cp+{�b�����~v�������!e!��;� �-��j��޽�<LO��ӍuY���f"Ya�9��Y
ᅹ�"��:-����\	�����s�����fN�����d��܌{�����5R��}�k���=�tm�c�+����<4	�����"S>x2���/�!(���rR���Pn�����������4���X��9t���6�7�����3�Ju��LT���觊���$鋊+6�	��N5�k�+��[���EsdhK;���]nˇ�<��ڟ�y��6�ii��R���_>���	N%7��uԅWrEz�gE��&�U���-l�)o	~f�2�%��*i�#�rB�.x+�����`KO�<��F�q��ܛ�uzW1�T߿��s��͟���u�Uhm��c�X��#t��jbz��ۇ4��~����8�r/���-���/t~<9zJ�a�$��TW��w,�Uͫq�{��綺��}��V��6�OX�]�Jp��*��g��9�XD�`�������<�iU:܈�6O#l;�*N�w��+�' ǽ�㬙~T� �l*I�\�NyBX˹!&8ޣ���g��J^9���~�b��Կ%غ1� �:�V#_!��X�����<s�0Wlľ5� �
|��2h��~1瓙�xK�N�����}�F=m��_w��˷v�D��*� F�a;��& ��o�nL2D������Zc�T���{k7_�a�����h�)̼����d�R����o�sC����Q�2��r��I%=I݋E�u�H�����8��N�='�W5�s,|����Ì�	�og�y�H���%?�M80`���e��I+������1�:R{ޟhLj|�=��Zd{mz�����Y��PS��I4����l��.)��U����(5y�$ܤo'�챫�^>���X�z��X𻶕��o�o���/���O��9���n�l-�9q{^�]s\��c4�U�ly�g�t=����:5� {	a�sI���̄roZ�{��0��OjP�9���j�Gf$��ճ��y��~z�o�o}I�� ���6�-��&&��:o��eU����z�_O� �}q�L���󭟟?���?����?t�1�,lՇ��p�i����{J8K��ne�<\gx�,��d=��lv>.��l6G�R���3�u��JVI��c���r�K�(vqz��/�;��ۋ�Z�&� ܏t���Ǳ��)
�?>fa�����\s0��E{~�A������\5��[��#Y�d���Ƌ�Ze h*GZ��2�]*c@����?g$.K$�j��o�b���#�kt��[[��d"���2�	�2�߸�أ��閴ħ$+��3��-��ع�+�%-��[�X�X�薇�vˮ�Qy�ɣj��ҩ��ӣ\��Ģ�������|
�q���z�D�Wa_
C���a�2�K�Ƭ8�;K-�z�^��Yv��K��rh�� \H�A��"�oӺ��/{yv#>�v��Jf[�Ī�
��Ӏ�Usz��v�wO������>V�T����+Qu�}�c>�ݚ�f,�|V(z��� �\�=���B��ͼ'ѻP�������]~r�����B0��_��	ɤY�Z߷- @a\#��b̛�`��ug;�#�e����K6P�XZ$�=gl�9�Wy�Zu?��,;U�A�-���5���F�+/��Ǩ�����f&��L&�3�F'��7�!p>@:8.��/\���
A�'zW Z:,o�>=�>_�p;�?Tר��熱'�n�Νk���b���%R�c�m)X{��1�;W��g�`����7{8�4H93��>"&�u�p{�������H���N>��}JԶ7}|(L�L0�F&b�ѤU��M����2������W����N�y4���t�}dB�3q�g^�[�؆]��:��Δ��尻������N��1t�%�q?�a���-�60Pl��-���)����asĬ����b��m{K��x�]���(k�%���qF�NC∼���C.\��$)/�ޓ#&��~6��22
֗ �l�e2[����ȂO]s�hٔ?�,^t�`>��L�0�^N���\�~>�c���I����EX��t���g�~sl�,�m/᭽��p�!��F�G����!� (f-\Ź	��*������f�)nZ���C�Yg�`�+j��9C����;���� ��a(c�PҴG�3��ʁ3��m��e���@������t�X�Pg��%5���%����Ń�~��%��  ��@�\��/����3"~t��EBu�49����E5֬�4���v]��&��z�\�T Yr�{��g=Ք5�}�\������#/��qd��N1>��6�q7׳�p#6B$��oeU���R�71	�4�]�,���j:'H�{Crh=��P�Y�.V� ��l��|LI�%OJ����5�eq���w;��$�y+�-�r�z�zλ���:�`�q�U5ԩ)�Z�o�)W@���u�GKP�t9�z�HA��E,W�0}�WO)�}G�hk����ʫ��6�K�ݚ�3[+�ȩ�o��j�J�)eS�M;SF��p�l[{��{,B�ƪ���'_g���
�+�	@��|�:��ݧ�K��+7�S�hn}Bp=���o�.܁���> �hH�����;�ӛ�r�n�jL����[:��b�w_�;Y���+�,Z��\Z](�,�×��DBp6�쟵�w�Ѭ��8�ys�ק�g��T;���?w���q���2^AP޹_$��"�W�3�4���M���{��{G�&RlP�����F���r_|�=�`	8����wVP���������40�K�}}QGl��-�<B���'���/	@=T�S�l����	�sy��l {�f:ro��X]f
�|����^ңJD���OZ���Mg�� �_g "Q��CPg{8a��z2d�B�?�v}�K�a2�7�4����?�A�U bYf#���痲�	��N�g_0�X���Iߏ:%�w�It���3|�/���o�(q����p"|؛]ƿ=���@m����;��-ա[S���yo��1�S���yNJʠ���B^���W�i��Wf.X ϩJ��hcQ9�ґ<��m5�J�#��T��ݛ��!��
�&@:Z%���+�BK��K6����l(�X��u�(ݝ������7b�ջ�P�g��Ͽ�x�@���c�䓴��?�o?G@¥��e��O6��#������U�Y��C�Xo�el���'t��Otiqa.���)8J_��l�#/v뺃�����g+c���g+���5�G*02�6��c�E�����)��Ap�5;�����ؔ��H��o�����Y&�=1��m�F���M�}�=G#��`b����׽�ϐ��q����2	q���v_�_��(��O���At�C�/��C2��W�k
�i�|/[6)�gf�:�z�;I�&�!��#��?b�/�������V��O�a( +��<*�ߠ�rz���9}w�e���m����k!���kYc띈�u���&~8�3]����g<y[ZQ���~�e�?!�o�p=�{JE���b>G4C��Mc��/��l��G�yR��#f�,%�����g"�Ďy�� 5�i��N��[k��W��#*��kNr�b���۩t]Zz���ݳ�
�V)���Wo�L��zK'�n�>��	��_k����%]8�E<�Xo��8+7D��n����jB�\V�'rRԖ��ZPԨag=gE���;cq���~6Y*�p��1�U���nބqM��+wZ�NC�j���HO�m�� Fz��]:4�a4����묇�5��dM�0R�W�1]b�4�T��v��:��r�k��z�T�Cu}S��h����VOyT̔��8�! J�ƽ�Bދ��I�:s��y;
"&���WiԳ|8v��-��[�!T�I${6^'��Q���[L�^�v��,7��|������S��F�&���2hO�U&m�6��@��Ĳ��AjT���A��j}��i��OP�|]g5=Z�}�^����:a��������{f���)� ��x����7]�a7Cj/���s�`Ȝ��'��%(�n{`�ˀiw}#Y�#񤄃�bS��J��]�f�2��a�u�Э��c5���\0r60&�?��{�?s�g��5Z���P2���4*���)x��j�z�WW(;}�mK�H>S;�dwd�q�4�rr���M��႟|cG�酉չwx��1e-������E� ��6��`���F_�x��g��]����o�GR�4e0�k���o}x���W{5�;��C�GF�:n���/�'���Rl�������j���r��a��`C)�B�/E�'~�G� ����Xi �湕���I�ܾ+�&�T�a�����@��>����e�����8����xz�Xz�Du��Fvl6�tY�J5(���_��RȰ�4ܪOp�S!�:r��M��ũ�5�H�n������v��2���.OuH����xn����Q�ϙ��w$E"�y�J���_EyU���Y��UDӎ�ED�;D	��ԍ�#�2����r�Djv�y��DOk��s��}(.vG�g��dP{��W�0�=�c�>��}v�C�a	i�+�uqp:j2M;�zɗ�&���J��,�)d�x����l�X�j�8ůn�����t|+��gSp𩘉Hw���M�a[�^���i��Pz�/ه�S�'�\s?k��N�#�3���٬qO�-��iӃ_��0f�B�]g��_����ʨO�����b.Y܎��
����A�pT`�qo�Ri�1b�����J��b�i�®MF�H������)6"�H�!�5*B$C�2zI	�#�|*q�LJ��4��~Z�O�2��qk���cj�8M3G�ӌ�����eg+��~:� K�X2筝M��bI\�QP�u�H�����LÌ���}�kxp��*���^�3����g�4w���w2�_��N���ḇ�	��Up$|�s�����bHBrm�����$2.c_@��򞣎4�~-���\ќ5i��w͗jPGTQ�0Fpd��)A����[#��g�.U�_8Bߛ(Eg���־��ģ�����LM�v�
pK�� �}i��Y#*���v�u��?�Y76t��̠g�R���{"KŨ�'�S���q��	����~/y��">M�`��F��,I��J�)y��Z i���k�wo`pl�,�vj���\�^9��#8T�����k�����(�3�r�V��N��<�`����#Z��ŅR]1�.�,@
���7�/�Q���"�	��Vv�L3sVQ毖s�r�o��w;��Fe������\�zj�(�VY���<�"zS�n��C��݋����!�+X�>��UU8(�^af*��%���M<��ޑY��0�.��jMW�)�=���c\�b]�f>g�1���+��>�<1�K�*�D���C����sO>k1(�w�M�E���$���-�r��f�Y���<�F�m�=�����	N.��u�J��c]�8�.�K��Xg����-_��&J_��SKS��*���Wv2�뫰?��1u�M�)\���Է]1"U6q�����(�sZC-�*礂п���g��/T�^{ƞ<��UË�f����?�"ס\���*�����eU��`�ΨBZ�����O	����;M�w��4�����!��o���çYQ�(�hǢ����?�a/��~�j�ߵ����j������cc�&�ʧF{R݄�{��b�mb	^C��Jխ�V��q�AUp;Gέ�^K3�(ݭ�z.�#����y���Pml��<y��Q�=���+z���MW}��Z��#���p�(ԯ���U�*"$��)�"�ԃo���O��Z����ݡ����~�M:dY9sȯ���2a_91K�!>��Z�s�q!��q7��Q�z�P��h����~O�DbWt�vX��K����/�}?|%���I!�ؽ��}�C����M?��!)T�0j{oRR�2>��N���Q�2��I������v��N/&T�)�GL�5�j���X�iA.�Y�)�Z��_i�7�"S+�U{�V;la��ޮ�c�3Bஂ�l��MOk�FA�e})�URC���1I�ۂ�q�OR�V�\/'���%��|��v��`��\E�V����	��Wm�*�i���v5�ef�Q�koC��j��h�_DF�cޖ�����+���S��)An#K��*�R�jiSF'�[�;�}6���³���9Xr��'wI�W���6dE^u-7IwH�k_�o��[+�D�n�c@��t����\TUr��e��_�ԓ3hF������w��	�ղ�h�45V7�I<"�]O�6vg�VP���_T�Yo�j{;i�)��AO�=��*�nE�t6Q�}�ۛ��q��$$�ZE���1��}ٗ�=-g��d׎PF����VNR���dO�Q���`6�(4���6�U C=��	����7�q[�E�-���=k;
/�4�nf�8Xd=���̬^�xW�iT��֦{�]R&L>�lUR(L�VS��Цk	 .���l�A�ʳ���>M��6�#�z��R�p�,�bE� �Iҵ���=�r<��I7D-T��s��X>z�MG�>j�j�O�+!W�0��5��.̝s�S��w�XG�Msp���ȝ̮3�k��j5ڽ/3��,N{�����7�ʏi��W�I�5�7s�:ǧ����=�|敏�,��]��L��~�S��;�h*�%�=�-K�"Yvh����ʿ�~�}ӥwh��޻�����_��S;�s���(�.$��w�854��Q�C����k���f���V6M��]���$�g�+��8xL�NFN����;�R1�4��=�Q_������=:<H�%��~�v�������x�c��Pݣă���hni]�|����+��=�|��BcJ�~����a~�5آ�4%R��2ZK�����R^[][�#��=�FE�������{���	�*�����_�Iy�׭�6��%�A\�Le)/a�9��)�/{w����%oR�)�	v�=�d�w���g:��Qj"@��:�O������D�UI��id�`��Xn���u e��@�����W�Wx�+�*�/@����g�B��Q7��7�y�W`ޓdƱ����c3;��蕘:� B�I{��~�~��޻�`��������X��l��˫�>x�Ζ�(\:�V�Se��pN��V��v���Uo���\�.^�yO�Ց��>-]M�$]�7zq&B��YK� W,��-��EmT�1�k������A���Z�88o�I.y�CxU�W0�5����z\k�|��.T��${�L��fC�r�� knQ�'T�5~����9TC��p� 6��.l,{�c� n�?���O��Y�E$�Y[��CA�J���%<�u�5�H+�>�����9,����7�Mޤ�z���f�����e�:�5��J8O|����2�=��kU� |6��j�XË��adn�~�����M�(�a���Pg��C���<D�� ����_J�U,�i�����f9<�5v+!�D���8������zV�[�k?�>�<S3�#��c;է�7��'�Z6C��$��u��M'I����(W]I�p�j�3%��R7웣d� ��_`�Li��|�6�sȶu� -�v��=��o��s�����˽h4�����_��j��t�!o\g��b�c_=�ö�D����}���9&9!P �Q�D���w���(�L+��׺�'�k�0�`��Z��8��(2�zB\©�2��)��Ga/K~;=���c� �A��~kdl�TT��kn@x���y���6I>8���)B��%3F�L�~���xAK�u�i��N�H�N�<��;�@5��~�q��?%�EX��0���ÿ�[�^����w/�D��`���J�Oz�����(����p��X��+�ȴ�toG�rT�6�%^�[R���?��oL�qe�rO��n�d#�7�K
�0�V���=�߱�	������q�KS��������0�-�tk����E ���+��&ʙd����ߓ�R� $f�ץn98�v�~+%q@,���U
d'���6�Y�����qw[B��%�+q�$��)�e���o�E0�c[���ń��R~-�5��*}k;�!v;j��ߋ#��D��3N��2�o/V?�V���8���0>��;�C{�."�6i<z�o_�MF��
&�0?e�u�&Z:{�e$�5g�K���S����Ie��O�Ͻ�<JZ4ISc-t� h�ROK�)�����M�K{*��yQEPH�K��d���s��i����g�x�&���k���r 7)1D�	1-ܤr�����N��}@�mQ��܄2R��ڻ��&�\o}�ߡ"Sk��z*c��w:�Q���=�ǵ��rV��#�D��B��ᕢ��f���ұ����Ϥ{��Tc�cYM��E{���x>??��5~�k��I|ff?��9����$�b�=�#!@,xzǖ&�*B/��V�������'Q��'=Q?{?�~����������h-{8ԩ����q�����q�K��un�斡���ESW���nC� ��{�f)�j-�� I�c
<���\�˵� l:�{95.��C���FD���:#μ�ߋ�G@H�ղ���'I{9{�PS��L ���K� �	P�:b�ݏ���(R����|si�K3~�յ�}`�zK_0�F�+�:�ޣ��b�R~-��މa��p��n��ޜ���V��aZ�����.��X��ҫV�����F3š|���%]�L�~E���B �֪Svg](��7F�ș4x�!y�~���� �KR��eﾯ$�=�#���e��Xk	s�R����� I�Ȱ�W���Q�§��Ԩ��� �(ة�����A`��t�o� ,+��-���E��$���ޫµm��m��ȼ����J��g����Qu�6VMR�����dH-���փ�������p(=o����~},7�_��`�7#���Dzr�ױ�����Jt��:3����M�UVdO��U��H���+}{H��g�]])��:�o5yW��n�Z���
~?�3���h�@���GX�յ�X|�_ą��M���k.�;�L��<�4����/�d�x+|�G9p�����LNu��%J����-U�
������ab�ELQ$^��G�	-�E����U.[����ɛ����(D���B�i�ߊż*Q��*x���RzA>����b�C~�u�y�f��?��>S���m�s/4+L�D�qRU��3�������ϬQ���e1/�E���	|Ƴ8��*<���~D/w���eumY��щ��ٷ�b����]k��͙�I�tnm�b�]����3�u��jjJ��P�хG���,{�ܛ5k���St����-Q�����%�kH�w�O;��!Y�be$�5w�ܷ^,>���ˈ5����un��O���.���b��}wc���N	�h}�[%��\4�����2v�La�U���lU��ն�^�G�O9,l�c����轹A�aN����B���f�I���6����1���������.'�3�L�ug��b��ř��6���*+��k�#�`�N���T������0�Ϟ�ƟJ���3}�����������L���PL����}�g<�	]�muϝ�Z��w>���ot׿�G ���?������ ���7ٱ��4���%$��8q��_z���;�c�w�?��{T֥�z�v)/Us�֍}H%��o�l��x�Ԯ��d���b���d�L�O�gB�Q���2���G���ņ^ʁ�o-�U
�����3��J�S�LQ��e�?w�gk��&���[z���o���� �f:X�$hy]�q�ӗ�g	�0�wFT�+�3;H�S���G��$����Q�w�"�б��Sj�3�NM�׍��n�&W6U,��U֨3�(����%���#�ǒzo/���Q����mp(z�+K�:�ܟ98�_Ӭo%3S���� *�R��V'&~mə�[�)L�1A���8+\��NY�.�9,RK�n{�v_���~��:�b�_`l<`ȤcP�b�dFUH��X��!/3Hf�v:l�p�=u�l����3��z�J�����Kvm��#���rgNe�މ�0�-oa�����#&����;�1�=CiZg�7-Gȓ����%w�����o��L�i�FP"O�Δkb�R>l&Etx�#�¹x0s���	r
_��X�M�S�~�U�G��zˆla������͔�)���IeD�\ pϛ���ޖ�����ΰ��H��g���ي�s]^���r���Kͱ�7��3��շ;9iZ���:<�]O�Ɂ��axY�5)r��ST����a�kh��.�,�u!<�D�d
��J]D��A��ڻ@魳��!E��7�%V'�l�_�{��������+>S���������i����c�8C'w�\�����/_x9R�⍌��n�xX����]��-���2v��� k�$��ML|�Lrxa�;?<`��j��?�2ÞƎ�hx���U����ͼ{��iM�ᑼ��P����
P-�.<�uBz+w��9���8~�۟��<�Sl0��Q�eB�7;��wT�Y�7�<<#*
VP��*EZ(:"�Q:���L�Pt��JQ� ��HB�t�AZBI�=$� $���� ��q�Y�;k�X�{_e_�w]���ݱaj�Q��%�'Iu���wi0b��a�+E�b��ĝ�_8/)3��7�h�Q�����Ѷ$�����sgGdz�0:���h�l��ώ�ZhM������f^���|�NQy�h����e�+�(�_��f�lV��[5/�������풬�nN�,�����ð;o��Qr�.��4�4��iΠzZ$i4���h�][u�'	�|[�j�ө�9:��Y�]NMu=����������P�;�D>��Zw]���?�z��m|Зc��*��v�����D�巍@�x���D�)ԩW����z��AS��H��d6`�q�F�x�5 ;͊l_��(Y�|=weԦ&KK�qY�����`����Y1����Ip���<�@�W>��N�D��>�,��3�o�+P�u���/��.�]ȥ44�}�Z���H&b��z+�m.�����L�Hw���v4��<9+�W�d�*E� �2�������]v�mE�F���Z{[�K�s<�� �K�n��|5�n����@Qo��-���f�U7�[rJ�Ԩ���$L��8}G1OqHFf��:-.Q^ѓ��?�?�"��,X$3�d��u덖��l��a����bn0�`lt��0��lx�:����������CX�x�&d��E����RH��%�!N�S8ʧ,%�j��x:$�:;�
���;{̬��ŧ�.��~����z'G��Z�W3�[C���Ӄ�^��l�|dظ��ʒ/D\�y4x��S����UO�g�J1@��j�9Z��2/>-��v�����%p�&��7H�#tRWɜݮ�;�K��T���gb�c7��������\���ni��Upi���^�
+Z��x�.�1�q��g9���ۄb��/�aĖ���2�WK�T��5����¦W�'@�qY�7��{����b�m�Đ�:��dY#���x!)he��瞇�e�g��0*G5T������:eF�+��Έx��.�;��7�<�f��*�Y�lwp��zZ��'�e0̊Y��Hv+�#��j5�������^���j�ZW�-]�$U�Zy$r�п���
Ez?c2�
^Jq%wr��=�Y���vr2�Ś� �ז�1��	s'h�-�͞����Ə	�s�4��V"'��p���/%������?�;��U��7��}�����]=��ld���C=�f�Kq���GZ��������;*�F�i��O�B����$ӡ�����!/��6����,�&���Е�>��&��o���\4Oa�9H�t',��77�,�~��]�rX�_bI�G	��X�4�(�e�����ӂ�6�Q�E#n�P/�>{ďt���M�w�~�E��:�l�t5��(։ڌV�ռ���{�z��-X�y1*7����?�oc�|��R�O���&_L��T�D4{&{'�\��;�T�R⺳�`���&�Q�6L̲ƶ.�b0%��-�İo��4�0h5����)�^>v�H�W��d،�Y����E�c�m�-�����.L������}rr�{(a�:\�Nq᷹8,G' �dbK����]��vw�j$�03-�8�m�N�Li)?�HQauvS��͓�<6�y���|�P���T��{��iC'@��_[Brs\,A�kbs��C�Rb�i� I��t|������LF���X�5�.܌ 9,��V�������nC;���7{�x�������(V�[n���|Bh������j��u��j�3K�ylol>�����kc5q�x���]yzS����n�ֱ�V�%��}+/V�� w�A����R=�8$Af�����t�,65[[fk�BR�̒��FPgQ�Eu� ���u	���(1w���-�c����¶��Q���o�%��i�-��I׌�!8��6��B��k�N?�����%i�jʒ�����%�'��6�'h5�Eɤ{��x&a��ȳ�Oh$狡Xu���;�J-�[�3�N�>��g"��	@��Q�K��c�m�6^"�1N����JR�&רȟ�T�pO̽P�A=�"
��k��2���w�0~O"j�{�A��9K{b�p�I�a�*��
�އLH���A\6~������6�N���.�T�b�B���JN�>/0�;W��8ӳ��v�i9�������7�0���r��;}ۡ����E��w���Kd�6���o��Ռ!��6���뽝A� 4�,�ɘ*�,��BP���cF�ي%�ʋ$^��<�E-
�Z�R�;Cm�R�c���
�p?���ufaH>���l;Xg��6y%_˄�׏x��A�Գ��JFZ��/�2�Ԅ�̓�b��'�5쨃�5;�LUh�3סg�#�H��ck�H�b��B�Q&bT]��NŹ�MX��V<KI%�%�o��4db��D<iݯydk�(P>�LnKY��;!"��4X6l�v9��	���G�A;����:�`�-6Ll|��;.1����oE!�yc�����=8��q��]���cA�ٻ���BK\Ѐ"�����n`h��V��	��S��\�9�*F�%-ĵ�.z[��N2Sy5���z�4(8�v�'�%R��_�N"��ǒE����5�	t�U�1!8�I��D?�~���NPLg�nyw�:�wڰ΋jB ]��R�aНB�`�q����F�I�aH(���|@դ!���5m%B1ld��Ψ��5�<9��<��lJ�]m&�m�6�3�^:{���P7��vʲNgؑ�eW���̳.����눌V9͍%jtT�+;#+�FԐ��yq��2�"z{<�,��e/��¸.�CIC����R��ؑ:( �W�F�p"��������B��"-�{�nkh��y��Zw��i|�v�PT]Y�� (�ejaC0{�qW,��zAX�k*��<�I_����֯uf��"i�&��S���0�;9v&�t�n��^�z��u��ۉ0�0FO��7W�s��#�.�u�"-fu��Go�
�2B����� Sˬ�5�u�����H��C����؛F�C8�ۡ��Ob�]�Z��)��R���803��������	���_��Nz�"m&����y���}65��*6���{�3�F�u�QØz�н~Qϯ��>��`�(����E)h^�����e0n�G�p�����i�&�lB9h+��;�έH����=������Hܛ˫�y�t|H1Nq�rWF�u��	��nL�r*+5�VG���,d�C��/�yb:[�x�1�r� A`���2x�{r���xs&CP.A�� n����a$��+�˦�N�JOp,*ǹ�,i�!�B���\���������V-�gp�PȌXߔ���I���`ހ�г�XB=3�Q�r>�a�h;jŸD�U������	�|�p%�$o h�+m�/vapS_�\:
��Q[�p	�e���6�x��4�1t�K@[��%@�L��n��@K"z&�+�i���/�=�mM���yxs4+C�-�]F��&D�z`�W���Έv�A��mt
1G���/�.�=\J��h�j5(��b���j`���}_K��]ص�Z5/W|���$q�:�
�`����m��V��Wc#�D�cZ��-��x.�ʩR��}��'%���l,���`g׎��������U���
�����?P̿H[�������ߔ�Z�~�5�P��e�k�I^�]z������I�v���Aʿ��~f���	R�v&wX�?�6)*X�&O����^\�&�{�����v�� ��B*���/C��?p�M��z"�	����q!�*X�猨p��R�[GX��Ϡ�s�6rz�ˀ�����bq�9�^p��ZeHF廵ۛ=p��;�v0��@�ءt����WŢ�>�n*�)����w^�����ڀ��M��u���2H<KXы�\��ݨ~:��P�6��ɄJC98�,�v��':�#�*��\A �(g���b��<�ٶ�ȧ+SCdM���s�)�x�Lb?V]EmL��>�|)�Lc���a<��2��
L�Q<���5~%�}�O��(�P?�������Y�:ٵ�6����@�}�Q�׆lf�K��u���EKRX�eJ5���0//ϭ�S���	-��	G�\H1�=�8h�c�5��U`��ow�E�j��,_k��'=�.|m�\���}Տ��g5�|�1,I�g[ɮC�Ê	wc����Z���J�&�6��i���RB��	�mm��|�Vf��kN�m@E5�ƞK�8H��Ϊ?+MTh�R��#��z�r��b�Ü.����WY��d�N㢂+��,M��DQ��>�vMsЦ�{����#>�u��?�WY�㘨G^"-�m���]+�ou7���S.O<�]�6�M%�BW�� \�k.�C9���������h�4�����r�E���ej#�#	��H�w6���V��/��!�� ���~�l����4?ҏ~�� ��LN��pB�m�QI�s9���b4`�^��E� ����n3�/_���k�R�r��zzg}�#m�,�!������'%B�����HB�� 2�h�M���8w��L�h��A#D�(���Cq�}c�w������&Bqy�����yx_9�w�������G��d�G=�.g�D���f�z�͕��fV��.�>*��w���\�>S>|)`z~��~&�7��L-a�]�����z+�C=g�����C�Y_��b��&��#�Ҏ�^���ŹŶz>���w���
�aה䩁[��u|(������-��鵅[�z0C��gk���<�F���I2�p����~���Ca'�;xxd�7]��1�ꗂ(ȿ^�}�[jw���9Д���"�;�<Z��q�k�k�B1�x0��1���l��4`�PC�����QF�o����=S���M�~�1B��d��C�)]��S[=�A��#� �_F�G�7��{��-�x�YU��X�<����#{d�'W?�Yu���a���{Wp���{���V��:��ьwR,e �$��mD���.t�}{K�(��?ź=,����s�� ����Ә��HO�KG�W��=>?:�y���x�g�Yw�h�T�~]GІg��������&�c�ѕ-6~T�x�q�U12z!����q����4������<�ժ����Q��o)����Z�ܷ�"�%��+�i���������e_U���>6f�W_֥�N���Q��.ķ+�wng��%Bm_����2�Ym�u��8�-3��kM�~��(�D�}�O�!�}t�孝�Z���)�c _��6��W���>j�.�S�Dj'�|���'}Ի��<��$��q��
�9Ӫ�1z�!L,Օ�����]��V���H ��E�ћw��{��Lz��(<ůORZO��O��)���w���+�8���$oس����U+
�r�^�S�D7�s�Y8�u��������wT��r#�Mk���*2�0��9�ڋ���un���P�T��P��o�z�������MM��{�(��~�����H�G�dɱ,׸���}�ȱ�b�*d��I���]��;�^@D��vO���~pujN1��]�B_5^��4�q�OYI-�~��k �!��I�U:e�v�ƒ��Q�\�>��w�]� ������9�Ԯ�`g�r䥳=
A	�M����gg�_p��r��O&x�9�X��g2"lz�mX��So�<
Q/Ʀ|2�dj���"І�E'���C~���+�	V�WPL#W)U�3Z���A~ rKʛ��Ƣ�PS�.KZ����C��[�f� �p$��I�ZF [��w�([����6�,P���WF2Y�� p�vQ�o_Z�nd/u�NR�¸�I�B�i�E-������)Z5���ɐ�������{���'�h�L4��/�"�y>ҷt�n���#����ƺN�Z��C~)2�m�^��6�OPڑm�� �%�|�\(��� X�n+��;z��Ф���ԟ��5�]�ҡ�Α5Ė~�p�k5F�s���w�o�)IV��W�C�]�g�-!@�)Ԍ�{�pۦ&`l�5.�.>4y/M�w衅\uNq��$�e���.{�? �����TQ����w�b��8�9yJ�/��#J���!�~��=�~9���(j��7וjd�!7t�h���&����Z��  �t��:-�sKj&?A�MS9:J���?7�`n�K�o��D'�`>�ԟ� 8/�.����E`����_�&7�0���h5������g��:�@�N:�n3��|�qz��BG� �����00;_�bJ�kq�åC�`%�l@�2ؙ�3�g���Qנ�n?%Y &e� L�Ia�t]�mfc�%�@��^K��- l91&��/����3�7]�4T��jK�z(�z }�t���t� e�<�+��M]�b^��,�)m�[x��>1D�Y�v���:(����m#Ȋt��ZY ୤���~'�,�c`�(*'u��k�ͤP�{Z�����2�[����(���G��٤H��x]L�(C)���^}-�s�̯3O�,v1���{�/>��%�k<�1T�U��X)[�,�.G T��N�P��,��Mho�����+D��W��XfD<���e�۰��y�`'R�K�	6��(��0p\0�����{  ��5}a�伝�!c77�v?X�V�}C@�XHt1��s]H��0���v�=�V��t2@x�^�:T45�W�Z!^�U��a2���
�?}St I����.1Ǧ�e����e����놀�f�ѥ���}�ȗZc���jZ 	�x,\	��=4�B��؄�~G ��;M ��0���LM��Q~�X��`a�m�y�hf����wޚU�r�̃H͔�$�k>�3ʳ��4��i����ʀÊ�E����)�[�gk w�'-J�>'������g��t?`o^r֎O��(V�ō��  �9m�[,���C�	$r�t;��k� ��9#[�z��Brl�M�1��j5���н���w9L*aV�Y]���E������KU>��h}�vwW�􎇺k&3&{j��.�W�И�͗���ǔ5!]_S&����&��hjG#��^��I�ۅy�Z�G��;^tKJ��P4@͡ڼ5�KR�	 F7�=��	�7W�L�>�la4�~����B3�eg������z�{屋*P�����^0�♸9ͪQ"��չ;_��)�D�Q�����K� h�' D΅"�d�G��� ������ő���'9��p��Y;M�e��P�IQN~A0֕����s"E�ʅ(�.^P�= <�F��.a�|�y�*6lcN/�˲�,~}X�Z��r�M�y�hgi�;@�g��w'n�����B��^��F�=�0K���;�-�PMe�yT�*)����pfV���maDanc���҄�6���+4�e��KGw̱�3Tp��kO
c����
t�M�]��ʴ��	�
d�/��x������m
Ta~c8mJnO{��η��v,nSY*�I�%ۖ�,F�q^,��~w���QM�~�K�
�T���T�@� �P�d,w VX�l0�x.|��a��P��22[�35��K���/��4S��xA�r���vyC�2<��X��"zV�zp��q7���}�#�Y·�?�i&���\���`4�]v;�E�	��̕"A�'Fc�vr��q3n`Xq�Z���(����⧆/O�_����]�������wsbH�vO���u��B������	du%�l�kh6'Y����V��-u��$�`�7��Xo�"A[Xi��d�o ��t_7΋F2>�A���6, c�r�hfE��fv{5M�c��Z�G���	���Rx��Ii����9�hjl����/���k̼Ak$Ԍ�L\�À�IN�L�Pm�xN��r�E��ȣ�F�_�!��w��$�B,3���̛�	U���Τ��U2��f�:W�!��n���P�+�(���������n�k"�� r�e�ʂ���EدXK�N+Kt\ߞ�n��Ҹ���v9�a'��3c&:�*�6�3�=պ�赭�fZy&����@	�:���jlP��������-�>�W�@x$�$�]{P�ڍ���QY��0}R�-�VH�����~Ҟ��W��YE�&�8�8ɹ�I�AS��&2�b��,Pj�<��O��dT)�u�-�w�,�[nJ�� �n�T$��/���c�P�Q>�<��ϯ���.h� 1tM��2�d��w@��5�k�8��h�Ch�jO;_����㺙�/��/;�&�V���>ˍ�W��K���w+�s�f������i��A���!%	�}S{]�o*bL}#+�sVΗ�Rc�W&��N
�7\y1*��K���Z�}=�^�#�M�Y����A1�}ۜ�T;�1�{�����\��<�#�^�x@�0���tK���sCA8����Ws�o|K�6xj�M��@�cKoל���IG|>����1�}�C�KlTKʡe�%S���$g�@m@�H����zLA�d,�|�>�Z�ԁdyA��1Kd�@�Z�R+y�l�	O���?�;�f�ܿ�T�s7#�CJ���A��*��9H���"�����s�����ԡ�(z4��&�y/��|N��<����n�/xd��9�F`�Mѥ@��(���x�0���:(7Gӷ��>��^����\~�Q��碛v��V�΂9���Ea���lR�Z�Ĩ8�$ A�M�9�o���ګ�VX
q'�@��ASO��7qc���&�<��$��g���2
�i�a"A)p����e�_9�0O�Z�{��ZM豂+	�&���������{�D��0�z�Y�ND�X�K+9�|t`�����C�/��o��rq`�N3�s��!!]��¨,B�,�/t�=3C�r�:��ۢ$h<	�Ƀ	����$nɆ���Ֆ��g�4FJ�Tޖ��t*Ϋ�����ˉYk�K-�� ��۔Э�MZ�5�5*�A[�z���yb�}�K�� �9��ëp�狴�E�p)�<�?��Z��E=�������`BlY㐊E�ح��aK4����-_8v4FB8��j.@���M�K���oJ��rzv Ԅz�`��IgՋ�r7��)Z�$P�����^���}��ܭ�w������D\�9]<�=�yzY�H%6*��XI0i�tqHB��I�jcm˝���.�w�������Ў:j,���k���q��{E�(AZ8�����A?�T�������ɝ��Ob�o�s8�x���Q�Nթ���?cx�>x\���xaT��=2"�v�Y�'��SD˫T�䰢�ReI9�K6�GVS0;�(_
�a�����dEO�?_�˖�'5\�veF�v�20J�>=�Q1;����iMd�v,��
��^�3���{@߸U}�{A�X�ߒ�U�Y�H��m�o��/�p��M��� �z%���޸f�ps}�Y��'��J9@�Kɋ�Ui��zW�|���&#ݜ����Wt��1 ��	��
#R(���i�(��!J�W׭t�Za]W���9��	�Χ��j�(Mh��f�<�g}0��|�1o��5�Gm����+�8�� &��.�<�p��!@���5ԌHW{���!|��!�0�L�6�yBL�c���!�/�T��^d0(�Ŭ�i�W��.��΃9�������"��'���C2o���J�1�-�[jC[�Ӄ�ea������dYN.�Gh�������)�'��;��k�b����W���C�ȥڙ2KEV'O��������Y��<���XB�TW^��6W�\�4�-��!���31R���琢
%S�1�)?��h^�N��(����Tx�U��.��KY�C��8��J�U���]��9#�Ī0�Q���K5��֦��%[�#"�1i���τS�L��>�BsS~'�0�Q܌�����@��F���D����9XKbg����Yė�1��hN��r����M?+�i܅ī�� ��cΓ OF˘>q�j;c�lx�Y����9�~8rJ�Rb,�0b��7'��Cwz�4K&8��}߁lf}P�o�����~��"����
t��/?�%K�I�C�Vל�&7�&�(���7{���a��e���L.u	p����KAW��\.*�-�[�r��d>����q��n�m]�am��L��"f�h��g�����A=��9(V�TR�Te�E�C�n�ԃӏ^r??v�N���wӇr���o��/�����.pu���Ts��:���th��#���!k��q^Dd�����v'cq��;a�u��]��O��.��n���`|�<���ӥ[{�.�q��zwi��%������,I �Pԯm�F�H�3@yn�#�����jG�P�r�'�]��\N�(̃ �?���lm�J^)_�J�6�<����i*��j��K�Ksy�r�(s'��u;&��pz���ki��R�RyKc�$�$�Dت�%�^����;���ȱ���-9�rP]d⍏�>k�Kz��߽�����,S�
�6�X���$�������4^��t�"VM1���G6L��m�{�ꈿ[vz�"֢GS�4
�۞��w��Ud�B�'%��iL"���:.ثQ
	��#<t��߅Y[�(2���xu�e��Dz� ��Ӎ0	O▌NC�;�S[8J�Z]�M�[Ec�('i����Ĝua���k�#����G<>2h[ZG��2�l�|�Of�;�!���c��R�"�B���]��i ��6M%	8�P%0�k�TD��_����Aw
�8���l�i�x������p׸��+�ޙT��.��>[�����&첚yr�\���nC�*��"(��p�H�`N��\��u�i�]Z`z\����!�6��;�+t�t�f�������Tn�~�$A�1H<M5��N���q��?��`@y�N�C���s�j ���.F�O8ٰ�a��ҹ�Ӡ]�ql�3�ο����9T�p���=������S�&/cI����ᚬ����9v���>M����5����=�Jb|(�wYMY�y�tn�r�(9�#H1�A��	���o�0UW���L����|D��<FVxd��r�a�yQ6�X1*�Q3���s��uQ ����0v�� ��$��.���d�Yb��xe�0�W��c�*{���(gW�F�/�ɰ�e1"b!签���Y༤+0T���a��j�zx�q�sUiq���jy� UI� x�M[.6"��5��]��t��p9��h����"O[��N#F��8����hf��]���Q���(T�e�`�Ĭ��Wcv����'X.�*�S��*�����1S�%l���%omjߌk��Q�4�����^�Mл>�震�U�k�Q��1�J��\�����jp)I]>� �7�nzz�Eͷ]E�)�H����Ļȅ�dB��E�IFT3�XD��vc,���T~��0q.^�&N_F?r�ې��Ww��ox&��W)}L�<�k�(�T����_Ff�;�f�/R�[ݥm�}~}bA�D5���ԛ��Kr5���
ȱ����̟�]�(nQɮp�B�y\��m�ƈ�q:�(�S��f`�I �g�Y�s�^n6���g�������WH��2v�n�I�^l�,��yĴ���고��f��a�BU�� ���J8��esq�qt���ǂ��������}�	v�Q�C+�7*�� ���}H��0��.*G��'%r`��B8E~����׽������]�g2���?d��l���|�� ��i��\~�p���I� O�8k9J�<p�t�)��8w��U ���%^{XԼq�UPͷ^YY4�E����M[Ϊ(3�z�|A5������IL��~�K�{��ȧH�� �����*�ٚͶ�M�W�{�5`(f���ڣ���ׁ�*ݝH���B�Ns����?�6qT&�����a#�	kS�������U�%�\�H��C��퀜���̠��k��>�)��@=e��V�����W�m�Fǈ�T��[ʇv9�Ԥ �W=�b#b��[>����Pg�7�+A~#�Ź�Qi�ZyH����i���e������%��e�$|T3-�`�o	��3b!�I:�s���ր�bF���4ʜ�|�ƱBa�}O?n�Y0���z���tT���bZ}�����0,���*���NPu����	����$�M��Vx(����m�vׅ�dI�?<')��n�݆{�#5>yu��Aqw�ecc��%(w���'��A86Z㔣@�롴ŭ챹t/({�G��X25�����i���T����������tϱ�̑��u��)��8��� �"
�N��މ��ݧSqq�%t�i�D�0�ڂ��`�_y�7ԓv��-�s>eM.��8(�zo�6��Y�IL�?������k�z�{�]�q��PY�z��e׉��^�q�����Ⱥ���yo�8`�_B>]ѩ
�=P���k�'�unp^���5\KS��=��t}��ړ¼k���݅ͮ	>Έ��K��H�I�w�,�q�����e�)�l�Ű�w`b����bϭ�+��g �T9��ݮ*A�M/
ɏ�%��7���KH/w;u��Q^T. T�z�yS�F��͈�w��?Z|CH�+��2S΁(��y�v�����7�[ٹ� �M�[�~�O��ޔ��M���\u���Č���[Q>���a�R=�5ӎ>�x�p���_�tx�ia�|��������!b5�_8ޕ����"���a���N�G߮r�Q�]�7U.��l%\���$?4�N_v�-6<Q8i|G�4h�TQc�8����Ս[�ֆ6�_z��3d>!;�>z<�Mz����2�%���v�=�Χ ���(��;�LD�L��h�R�p���� ���*��"��/or���b����:��UR�����Z��O���w����R����wew�:oUy8���sC��b�,O�|�+֘���Z7�a�<я��>N�����|T��y���ap&E�1�BI�~��,���a6ÍU/Z�s�Q���n�u��
�|���:7P�]��1{M��1T�=/Q+���_��CZ'�Y^�>�?0"���w�4�O�xJ藮0λ����k�K�1������-��T�Ae�F�GFĳ�ˍ��&:5����v��[gg���Ptڷ�;�������}�)�4�hD��:�8d���'vA���}��Ȓ#�,�7�!?��GG��w�@�`Z�ŵۺ�!:���k2���m�����v�_�3���,���V_{��t�{VҲ%h�p��Ǵ�O"�c�.���cF� �=��mIE�޸k�O�ɁR�
�@|�)����G�0�x�K�&�]c���S��D7�2��N�����Tu�����5�sַ����&}n�/�P��"I��>��J��L��>s�+�X~RK�]Vë���>�y}G��G����q%Ճk���p����9{���Y����K�ǃLJ���x���㞮���C��S�[�$B�;�'�sc�ϟ������̧Ge/����t�E��9�{���1��g��EOU�ܺu��W��؎�\Z}
U�On�T:Aذ�����ɨ��r�c���������;4x��?���h_��Y�2����. ˜?f�^l�VsmI��ۡ� ��;�?e��j��gm�����,�"Nk�ZC�㖹�B������6��0W�?S�g��L�>�� &}�\-7�����(����7c��;m7Z�!����M�#E�T���$@-dg�7dn|�K7��#N���q�������g̕��v�'��d��Qg����������Ñ�e�Ѻ�.��r�H=t䟢E���м#���q��D���ŕ�.Zs�׏��.�gUm�?��;)x���骧ǿ�PС�'��������o<��:�y|}
��v��1�ŘU�5���]���N� ��$� �"���H��r�a5��ǫ�^/}��:r�,}.�.tX �bP��Q6��"�Z�Ǟ��O��V��kՁ#|@���q� ��G�1~����3���S�����~���J�8g�w��{Τ����H���t���o���1R�}bf��7��*�H�-��k(=�#�>�\����R���H�������]�,u-�P�;��Nj9����v}{�R�=���:-�_C��^39����D��^����?�rT93����
���S<���zn����#y��[m�4(�A�3�DsH�@P�#C��O4gG��N`\!f�Wӟ��b8Q"#�"�e�ؗ6�Y\�������1k�i�_��oH����6Iќ�\y��SK��':w����>�*H� VL�7�,cq��?�ų�p]Ra��D��xi��Y������_u�b��~���#�t�r���Ma	�\����n��^���*hM.�=��0,�W440�%J�x��;1��-Wy���<m�����j�|C��E���l���\��:������wzݍ*=,"ҵSٺ�v�Һ��W,&xb���A9��k��c�Q֣��S�S���	A �<u�XW}�;�����X���Ek��ȴ�K��S�TV���'e_"��/�R˵o[�C�+�pAs�gba�x��]�/%��!c��^\ǌ'Q矸�i̜���!���=RSU\���2�R�\�9�T>���ߞ�Z���a^MC����j���>a�Ã�ŭA�'3��3L�򀴓�߄�ٸW1da�O�_���F�����3P��_�~u���R8ak��ZWnm&;�.�w����X�����Y_)LP��	��k�{e�nH���&�B����xJ���T�~P�#��q��S�S�<m�5i�qv$��ק���Պ�PH�J���sc���U�$��%�5��y�:�^��K�|*��7*�����ֲ�g�JK]��v+x*5�вl-	Gt��Uש��*��K�e�L������r�]w
1R1*��?�yb$vp8 *	u��5�	�L��(	bF����P�."��k&?N�4<q"�2�w�D��ͮR�$�w���ʳ#л� Cv��~)���d�جy vj���ņ�`V��K_Oj=q���}��M;��粔��eP��l�bTds�Z4;f���9���6�h�;S�^�5��X?'�N�IE\H�HϪv�s����4޺�cM�{V�:�q=�
�O��r�>���g�B�B=Y5�#)������n�4	&� e���UW�+sLn{$��v~h��Z�/��(�ᳶb�,����3H	�<�)�.�{��e�����M�iZ����$�j"ً����ol<�Z�%\�����%�_�����GC�NL��2T��(&�|(aG�[�V����;�����E�D��]��@� H��u�ʱ+V�	�|��t-+�����[[ۜ�:����y�E�F3?ٍK-2]E�Ҽ�#�̾��s6��6��DIY/Χ��o�]Ag%��	�(��5�T�Z�+V;��˚{�X׀��b�c��T/�RH0�t��˅9�+��dm+�@�46Z��ц�Hz��h�V��2�9;=7=����T�F}�JLd�ɨ�P{����M�+2�j�dw&2q�ڼ�ZS2��@��M9�LX�
��9�����!u��Ov���j�%�sM*����@=��Ft�fB��X�t��6�����2R\�L�a�_yl���__"�K��nm_c$D;���(�B��,�i�rM2r-����ދys�gQB�H�r��b�JG��,ia�:�Q��mw��]��㥐������G�� ���� F����k%	�ф�}���0���P�W8|c_� (��eI"�0npL@�吵(Y�^��m�7ܝqY�YK��hF�΀���S�5������%ӄ��p�S}%��������0aQ�3*������%c������oCI�и�����tw�b׸�Ԉ��d�y���Z�aD��&O�&�#��Vzn�T�F�FT�-h���a��9�ξD�͟��Sw	����үq�icu�_ iŞ!WC��Z뷩�3�r@^8��R���q�[��?n���|��P�/L|`/�����bj�^%ڜC]q�
nl����jM�VoG������-l҂t�H�ͶO�_'<�cj�F6_��T��珮s5��.��A�!]��J��m������̨+iKJ��MO\~y_Y��"!���kTZV�zZjj��5}!%曇�w�9k��J}�ۑ�t�0�j�WU�\��I�R�Ҡ�K���:�2݆��$���^ʭ����y��8.���u:[@�f��p�׬��]�F��t���s}��n;���p�<���H����6^k
�>
<���sg�/��ϵ��Hy��4q�R�&�♬O\�a�UsZ��X�O���T�D�A�#0Gq�S�F��Ћ��=�L.��8�L�VY���Lζ횞�@�{5_�FFa#7u���chSO�V��>����w w"�,NF��,j��??`�
Z��+;51�I���/o���:�v�����{P��\�n��9�62��~2��{	"�;�oPh��)�[�C�����H�Z�!m`�G<�uL:�����Fc���ɡ����ɩ�_�)e� Qm��D��ʡ"p���X:|��5��
�!QߙQ��(!>���&�Q�gQs����4���	���H�㢺���۾��A��s�>&�_`<O��(B;�i��ݡ�<�51�I��W��=�ڎk]Ea'0n&$km�#���Օ��Aas#��˽\�2deH���X�I����:9�^�֠���UV?c)�;�"�`�5.�+�][����-x)�]۹������y.���L,D~+L�O����C��.۝E��@R�o�Y��7>A!�5��*R�((���Cٗ�L�� �k*��I�>�-C`n�酋�0��v@�	��R�����1+}s�G3O�Lt�7ȹ�4M뜷i�J�����{G5��}�x8����"�
(M����T�JB�5B�MS�J��"5��IUj�5�P�IHB��.�>[e�q�_w|�{�x�p8�bΧͧ���5�2�+��Lhka�G�t}Z.E�B��r�iw:�S0,�Hs3�� �������z+���y~�2ݪ�ńЛ��?V1o	�k�����֙���h8���8������>`B�})��H.�L"%��sS�l���U��}̪����k+�V���L��<����6�k!��|���߰��˅�=$ο\�k�Qf����$�J��4[���~ԟ8��Q�~2�/=�U�B�I��/�E̩�����!�LA�:)�~�-��% ��$�q�i?M-���iU9���S�ʑbb�1��'�#�2l uFś��K�{��K]N��H������4!��i���rq�-ȯ͆d�����^��0t=����p~K)�W B1\
q�t����'�>#�z�(H@ҏ/-�a�X��㆜c(����]�u�'���$�d�l����A@O�D�!�ȳ�)P�ӳDw��O�
4k I^��mј���Ǘ�(�1�ڏ���H(�d����'�������c;�r/"U��Z��׮ȃb����9��u,3�Ғ�N�pb��`"B�%B.!(q��h�i�%!����O=�q��P�P�#�^�}/���@}`��F�bM��8�*�s���Hi��e���N-qT�v�ke.5�y|H�{���見�4�G�};v�`�c�Y�Xh�BJ6B�p�;
�>a�	&?׳kP�=(UI�+�뫐���<�V><��\G�q딬�Ʋk5�nT�E��^)�e�|�9L88��q{ލ���}~B�̫M��Ő����i�}$T�\�0ݐ��/�0�l�M����Kopu}�\��f\�%��e�J�/�d��!����Я�,7:�!$"��nD�'��Y���>�*���Aγ���{�T�A*FL�@��x@C��-������Đ��N_/3Bd!�F��8 �0�ϩ׷�is�&�Gw��,>�����k�1��K-��{��r^��0��l��Y���2��g��|�t��������w$s�~�%�׫'�>w%���?椈�技�O��\����v�9Un%ÅC�7�=m����.]��l�1��W���6rM`h�( z��XQn�j�JM킑5i7<�	�$xw�&���.F��Џ$V��5�y
0�Do�j��}P��ĺ�J���IXcJ��n:N+��B�OTx-4�r�3VD�>1��J��n�Cm�Ł�X��*݄ �+i�,���X�b��1&S�wj�u� }�H̙=���o�����,�op�kk/=�x,U{�r���u<�	�= ��Z�^���4B�zRX��tE�*{ֹ�־�jKdAp2?đ���Voϰx�X�{e��y�����X���Hg.\���2��rc��GL�kx����)��Z�^b�_�M}k���,�RW�@����w$I�w���:
��J<F����%��HV��6���Q�:���A�쯭Sq)Pbi��@3_:`�Ur����K�)�ɘ�^ݖ���DK�VH9JO��h�q"@�5�QFU�N��>����Ϳ��&w<r�vV�T�D��%�D�قFҧ�\�h��o���������,AZ"��qM����g���M��mv)]Ũ|��ϋ�>����a.�����ģ*X�rl0��1�=K�D:�t�od&8�CFhq���V��GS2�)�!$ޟU��w���-�m��V%Pov�=!��g۾�=�Sb�p�u[��e�[� �I���E��Ab:�F�Jw�������ĬI���ӆ+x �ĵ��UNv��3����k3�l�I�)ʜ�;F��P�lEhåX~��+�h'� ە?�w|�X�j���
m��2o�K��}�|k)��=�/'�Ww8���/�`9��i���W��[q���5#�? 9��: OL�Ǥ~#�:"Z��J��L����鍫�J]����M\D�m�[�þ������a�
���ɛpfs"V��{�[�!B�G�q�i�!� �{�)l7��vc��%�)����I�__�[[}�m|)r_ze׹W��F=�p�����Bׅ�!��<����a�|Jc��`�͗%�ʼ�߫wWY�mm�)
� "�-����H!�v�	lS~�Ǘ��[�!%����5��ƥ���T%C��+�؟�"u,v���Щ ���C�!�G���ī���Xv=�,R���aP�D�����A�	
/G�=�)|ֿ���.�v��e���~h��  ��P�+����bto�f����߂�j�ku\S�gT{K�v�nv�C�v^`5U�1�V�D��zX�!��EW?�FEh
-�E���\&Ѿ_^�&Ͼ��	}�?ɾ������<���D�<JR�z�+.;��k��m��E�/V�5����p
���˯/���@� ���%�ǜ�Z	�e��a��+���.����? gM����/ u�=��s�� ����4����������Ə�_�J��M?�F⺭$DS��'��ѡC�ſ��M���㛳�e�U	g2
z�h�K�g�� ����n�\���Wg����;cdd��XM�u�a�z�F�ֱ�o�9�Y9�ԡ��2J|4&ꎎPI�?��Cq@aD�7 ��������Եoov5����y�YͲ�&�)zW�LW��p~���A��g}�?;�7�	e��ubK��t3�ht!�r�oh �d���Θkq+��?�zY;�UZ��&��%,l�g�5's8�b�Qߘ���3:���"mʭ��oQ ��ugߑ��X�b
�߹i�����<�ϥ(�E)�ͻ�Y���F0��1~U{êaB	e���� @󜫋�cJ��Jl`vW]����X)W�M�moۚ���Ur[��Іq�������7!������.��k����'�� ���r�sHX_�?; `�K���I>��ߞ�I~�w|4f3Af�С���3t7�H?�������Z�-tJU^���:%
u�I;`�eZ�ǘ�13k�5�!�-Z�������B���GI�^{;�Z���e`5�
r����~�e��Y�2}�|��r`樯҄�孬\�Ǒs�su<�RTT���4h���~î<1
a�X'u��Zt0��گy1��%�s\5���Dw� s%F%�}�����,_���򾾸��r������:Q�U��\v�	?�zm(�s��m�Lze�� ��<�Y�l$�09N<�rZvA�򓚧&�mr	�]op����ؖ����),������3G{��u^�Ǿ#ߒ�j�Ȉ�(�UءWO�ϟ�ZިU�Z���,���s����d�s1��G����3��~j^dR������H�٩�:���3$ރ��9^��3 ��^�;v�vN�d��*��|ǛB$ħ��V@,9g�vf�ZP���+jNx������;9V�>�k����B�7�w�(bC� �L/	�c��f��D!��98Ny��!Hʢ_�C�s�t�@5rl\�26JU�$��`c��C���G�d���f&5�`1&��9��� �(hw����@���P*lnh{�J��vz9̫%У����K���������T������Vf*�hY���]�7OZ���Qt��IØ��G�;�vƈ�m`�ȷ�7|=:���/�My������(w�jώ�6�: ��`�6=q����g�����v��[�9_<Ro2Q�*v4s�
�e-��[Ԏ��Gk��K��w�(A�G�||�d�<���6ޏ��T0��iZS�7l�����t#i�s㾵�I�9Tb�qG��[�|M�N�p�~*׹�����kY�p�p5FК��#��xj&*�z��~Y�Lv�ȍ�铐�ҳ�!P�B�k�fZ�k�`� �a*T�E� Ewٔ�f���s.�P"�t�
�����������%��qG�j�;�'&q��a��^	2���TR��I @���m7�M�W۞
�`�wA��ϱe�X�g#|���ے+�%^+���KqF�@�ʳԒ������w?�ׄ��{پ�z�>w�ԏ���'j��C����;�B@Q�J׃͎<Y��P��r�}��{�����ψ��7�B�����qɧ~a�@�R��m� �羠��.9��6���v[���h�C�P��_��0��"�M�{�e*#/�W�e��
k1��Rz��y�E�G�S���p�(�Y��x,CIK���!���.�]߫�o�|�3 &7�f#�SD�Wm��ܶ��E!F����� �K�il���#9��|�n�f,�N���s�����y~^���->k⬍����u�o���A���ͯX�*A^Xo�L%�,������%y����:-�F0�F�3oH��X ގu��q���e�Q����O��������HD��_) ��>�X�}�aO����3{�ݘ�E=�4��0�T;�`��y��o�YՃP����è�7vf��^9����5m��i$�?����`�Vj���z�@%a��=�c����Fq�:[?�2�m�x[s]�}����[����
7�����D!=�oب�^+%���=B-Wעӫ�쇫$-"�\	�Jb��1�o��0�1߶W�z	b�q�f��G[�1f��i(�s'I�/}��� Yp���j� gnÓZ�<wG%���X��+/��I��'��bv�H�����y�ԁu�:�$��硙��/}��Dݝ�ӍeN;�WFi��D�!}�@.UA}/�Q�_��{_��������� ��Q����8��m����b��Dַ8��M�Z4ql�o��.��-�����Ę���sM�����՗,3��{;�n�W.U��ۑ�%����"M��H`F�4�&׿m����r(JP�PK�� 8�X:�ߠ���m�v��Ό �� w�"��Z9'3(p�sW1�`x_A��z�z�z]�@��v�k��f7�����Ef�ʚ�^S:��8*�?%~0h&��eos�d4�=�A���5GOmKXT~���Z�VJ�ɍ�u]��cq��v?ہ��`�(��@g��ɯ]�H��8P���C�}{*|�ѹ�(u�?!l���R�K��3���ȁ��L*w?�6�<\�����ԓ�'P�1$��l��5&�a=H�XmPW�o{v6�66���g\0dаj�ݬ�PCŃK��j���' ]3�c5�}�Pe�����Wt�1<���F���p�=y�x�´�ka�����l߷T_r�Ha
��r<h�f��x�3㿙/�M܇�@9�vV�f�n�%��:����>gl��xAc�����Q=ح21s�-F䚀jy�U7!͏ˍ���5����P2oP�X�w5q_֢ɞ!!�(3�	�\��|�,#F�W���t���0٭)�mI�k�t�o�",�aDLU|z�����1��¹F���Ċ�w岲�E	��9��{�IdP�( �GS3�V.`�X�����>leD֤\IІg���e�4X�������\LZ��e<F�7�c��7
f݅�,4K�btg�Z�|p�e�a�ֻ�tA�~�3���N�������7��q8:i��Aa*vS_���t\OO
�,.z��tg���
��2��f����;%����n ���pۿ��3���	�mD��׃Z&�*��%�ԛ�a�)̐��EKgB�J~yAy�%��
���w~B�$]��N z�e���M�x�7L0���P.$�sI�H�Ȍ���B�D��[k��6�x��U�/�|i�X�E��0����r���@t[��|+� ?�#����&��Z�yZ�ȨE�fx�.f���n��`7E�ѱo�� `&T(C�fg-Bls=[��nvx��w]�|n���d`�@��xbl����~E��u�r�M(,V)Nk�����a���a,�5���,7o�!��E;�����c���&�Ҫ2kX<�G��X�/qR�͇{-K�*�E�Y�2^��f���@ݔ"O��cW>�r$�h7�{|n��R|+"MŠ��w��'�Dyz��L�\����^��U���"�p�"z�a��9��ӳda�s��m���#Q������78�؍�@��{a{����\A�p#�=�<u�SKQ]�:����v�����F����0�]�]��F{�����t������A�z�(w�i9jj��?x�p�yY�]�~�b�nL��ꋷ�����|�s�5��Uܱ�5�w,�8��`�x "� 6����O��<�]��f�`�ePa�֛gP��k%u�7�����'�@�5��.��rE�De0�������`��X1�#���KkK�d���U��N�*�՝f_R�蒁nvc�1S�Q�+/�6IǷ�~���ߠ>��#��O�������v�E��{ZH�,7�1�s����|�mt�:���!�(?�%��U��lpe��V+��S�I�ΐF�A�=ʱ��o�6j?�O��~,���mbu�s�W���+$հ�JQ�ff��'���|;{5�ّj,w��s�f	�����G��ט�qN�Ǉj�v��.8��<B�|�y �����t�K����jnv���U�� v2��z�z����Kx���i.|�Whm�.�����rFv2L���4x��a��N2�!�8�Q���Χj��#��u>U f�Y�N��+,%O`�sJ��Ŀm�,��6v��")Ö�g�'���`��}�KM�^" |
����b_ly�困1R;,��V��Wk���<�a�D��᠊T���V:&(ѣ�������d���1VD=^c1��ȣ�fKH��E� ��X�JFVڔU~ed��En��8r.DH������B�� L��$��خԿeV_��h?�E�ت�[Z�2go��n$�L��b�$+3���4�[�2[�;�� 2��"�K�Ap��%Խ�b�l��ÆGv�C�U�]�A���U��@�Z]��ӔD�����pWt�5���j*J�6GL��aZ|���R�ĸrI�w�.	|d{���G�JKyI�Fm.�\�b^�J���ռ� m����W����4��	����o�וP&D]9�h��h�~�޽����0�L�
Y���n�2�uwB؝���u9B����2fI���b�x���8���%��B�ƌ���*d7���z�H@��C�� � �M}������i�x*}/�*X�W�0o�*>�:�C�b����Q�{��(��	�XF�d�_��ٳz�jя�2:�^�b�N�x�n�NeYAU�~2+����z�c�`3���d�{�L��դM�a΀-����f|�2���yij���M���I�sI�
>^ݾ�a~��Tu���`�ࠥT*'��ϠL/����Ȉ:��y^�P���ያ�������ݟl�?̒�E�>�צEVy<�^�VGe�)w��/v?���0����	�M@p{��PW#�Ƅ4�9�TO�t�;�Dq9��{��ñc�����v�ug��*7Zڀ��*���<���IV�nq�be��;�ߝݬ$��y[�d��lT%���Ae��W}�ׄ��f���]�<G-:}�e+�����A��,��f�$N��QK0ǭ��C�3#@}&8���~��´�5Ş\� ��ڃJ@�(?Ѓ��_��p��"LBc� �&yh���qfpCQ	�C ���F��P�{�xk�,��\&�
B�2�N�cJ䫎��M�-��x!�)�P�i����E�C���[>H��^��j8���"������Cc��&���yr�?Pm��[�gH]���a��!3pąBN  �E�H�?H����������S̠���s:ˆ�UX���J�~�6��|nJ^�=�z�PEQ5�a���&vw���0�|��z%�
��p���&t���r��am��ܚ�J�iGγ�
1`�j�!�T��j0����#�\��o�Z�!�vD�>?���Jry��kY
�4@XwD{��6��g��-���>�i7ZO�+?HM�������������Y7J�F�Tuv��0�҅x T��-l,|�Nb���؄�����|ܵ��1P���+*������_�N���[KW�X��/"7la'�%hh�}-`��.�С�\�x[u��.j��`��*�~�ldɖ�wp05ȭ�9��[��"�N�Nu:�e���ݕ��=�6(U;������5��.��B��N� Ƈ+��X|���ee�8�
F�����.��<kNRG^���"�|�m���6�I�>���%�l����T���k���g�d��OI�ɇKK���I��o{s@�G�]$����-������u�rӲ#���j"����_f�C�9�
$�_**���o@ɺ��+	�ꂔ�v��I�g��u��oP�2��(�;F�%lxmϖj�a�v�78��1�,�E�����d�����.D�4*H�m�Ԁ��K��s�c#��*a��)�<�Iɢ���B�,�.���͐!F����5gB�Kx��-��s�ZZ�Z4�K����R⹊��\�L�X^�7�PFA�V�''USY��VRp�՛����R�������{S;���w�[v��	8o4�8�	�8�L��g���2�{��:袌o�M�E�a�TH��d������%�5o���r�,�7��7=\O��PFC-�Jb�t��\�NC�e�`�/��>��M�HiL$]vf���p	�={�T�2�b�8�)9E�+2w��.���"��ē��>6q�C�=���59̐��7/�����Z�88���v���C.�N�:y�����VwN��9y6����2�O���_���2�q��#�R]?����ڙK��u�������-4�k,c6q�cN�Q�;���k�Bh�`�:�	Q��8n���JO#/���ɧ��G�Pr����=b�����`?������P}i!��m/m+X���vN��|����]qU����.�L�'T/˜R-�N�����p"�u��9�S:�A)�#I��9J����]�7 rE�����!ɧ�
U}F�R���"瞛S�3���!ԇ��A8���.Fh���Ј��;�9�T_��XN8��\����,��ꤖ��$�eI�J���`���؟e��[<��O��)��eh�m��e*#�\���J-�ow\6���@O0{k7�_�Z��{�
j��o)"�'Ѵ�?�#��r�( ����:��ȤW�0o{��DNQ(!|y�{~)�9PhB�C�,}Xp+��0cQ����ܱ`���X�цH�jNHSa;1�6V%��6k�\�0ޚ��0#/'L��_
O~�k�y�+��M�� r�˂��-�۔�ڼ[+��@>X��be�E1x�{����s�@�O�?��m����U�:<� ���h����24��[���I�q�;�c�ߐ��He�>�c��J�E���ꇵ}9�ǹ���e�HS�e�)'�W�`��a!����Ӣ6�`�ߵ6��!���2���'m��!����u mf%M��&|6����˛ o�r#�qrBE�!�u�� �j-����/|t��q��׎����a���$y|��BW�n����v�����;J�\�@�v�i����{������]S�R��X��K����s�Boȿ�*��p�,�hP����c7LDP$�����\���:V�-MPK�F��x��Ѓ��;��^�G���o��Ei�� '����CKXr�Z��0��p�����`"pb<�HuK��`�a:�5�fT�p�d1��wU'���U�8|
l:��;!�!��'����o�����2�_���1}���wH9�+�����fnBwA�v��VE������+Ayjv�D"�<i�4�З)��X�.�`���y&ݖ��Nz~����=܀�#r����q-[}���[=.�	���	ư����8	�~��tvH��30��m�jy�R����ك����Z����.�4����"g�Y���d���&��-��Vğ��li��$��S,� )�,^�.�eG���
q���3`�*�x�,7�c�"' ��@�k� NZ�.�<~`*��W�Z)�Li<H���܇6��MB��%�J�s������������,D�>��-��I��Ʒ������K	5o�k�+�:�I����sKo�Q�3m���z�F �����>Je��||k�����Q�E����\�E�h�Le�z�a�M��2,Ë�ɳ��: ��t��п1 P����0�œ����+���9��{�SAF^"@�t 
=���AV�� PF��ȏ���K�X���1�3Z�q���obqg�.�5,�".YU���^H���
0���O���e̹L��V�mu6�-��&�Y����f���NM�_.�?-Ks��W�\��,�����9e��$d5t�Il/lxb��3��Z�>/�<��.�����տl�ff�n��S~��}v��Gå�9fN�;�2F�'ࢌ��,_�[}J�<�)�Ex��PT��1�9��]G���H�|�9𧞳zx�?�B+Gw�ɡ#;��:�Ò�V���l�s�k��~�oN|�ҁ$��uGȋ���cdŅ���$v���B:���J�|���*���j�[,�^�fߺ��vL��=�i���1?���ඵ��>s	L��E���������=�ҍ�G��a���!��2,�7\�#��^z4�7�`�+D��6�"���� ���#��23�}��(���0L�c�/I��ga22���w�?�-�~��G��߃'����c��1�Ӽ}�f��뎙��}�o(3�[������:A�!d �#�,s�+���jy�q�������.�Y�R�PMPJM�3�j~��6��u)v��~��?��IBw���۞�9��]���7��)!��z�]I9
�WF0�g~���� �ph麱� ��l Ud�ų���D����S������e����a��-7�m8:��Ǽ�R���&Fs���Z��i3��ܠ��&�ԓ�\�g�zճƲp�v��n��E?>�Q!?1��3}�ApSg�� 7Y7j�8���Ym"��9�1�f���1(�Y�{�c���IG�]�GyI9��FN1�b+">�m�J�i�����G6\y<�w�x����|7�16f�]bҧ �?����� �sb�o9<�G�Y�m��(�Y���Gx�<��0?���~w�J$�u���۾?���� �+O�|�-��
�^ѣ3��f�M �[����3ԦN�(���������8|����_uj�Y���b�B��8�-\Q�wM��ZNԉYd�f��`���Oc��C�R3�o��9��P�34� L�NL{��1��N���˧SF�r0�jS����Z�f�Q	1J����ӤY��)f�z_�jd�q833�[�q�X�#'M�Kl�ع�/�y3Nk#:;��\&�M
���6�6?z��G�o�I;�Ƅ�ό �Ԭ����u8E����}̉��-�I������V����^h'�i�AĒ�n2�C���m�;�y��~�jn�O̒~���s��g<�s�ɢ9T)>��J5�g~��r.�r£^��\0�t�Z��E��r_w��-�2�(NPW��Ihϲ���-�,��Z����-g�
]����@]����>݉f`��D��oc�H�٭�s$2}�).�o�\_����C�����E����1�z��P�;���WO��M;0�̶
 p�e>`�*T���,R5̔8��s�XT��3����A���A��?��� �~�s;b��p�6�!��4+����V��9pG �Q3��h�:ԧ*����eD���412���?Vu/]��6r:�BW3�/�~o�` s� ĸ@�f��(�L����8�lՑ��U�1m��6[[?	ׯg81α=C[�=��瀜tڃ����rN�����o	$�]���|gX�QT��ۙ�*+g���9π��ׁ�=���g���/v2��}U	�y�|@������M��:v���?���y�����S� ֤S�����4��"���5�6�sN%��Gs�y�6��O����n���V�|9N�����7��TT�t�����7�F���%���V��������xEsV����z$ne�L0q������@�i�U��9W������^ssv.�?���H���V�9�B��h�C:n�����=5�,^7�n'���>H�>�V�U�_sd�W@���E�\Wqk�9��jh��7{������aq�g���#�e<-�x�#������;��5@�@���l_r�O������s6#�[	LΗu{oi5���W>��S�/#�P�G:C���)=P印{*c�`O�b��������+9DgC��;�HX��q�e;\�����=��a�9���\t��ZC�!l)c�_�K��^���<����V��Ay����}�\���05��F�*{�x��3���]�](���27
�_�lgvL
���,.�y�
��>R.x��5k] B���(i/y��B���7�T�J�T���E�X�D�X2z�O���
��I�5�I�7{���Żo��z1��A�sa�<A�-sH���d��!2%�}�L,X`�uż��{��q�����a����AAT��ƅ6���b���<Y�Ve�WJ)5��>G=�6��0�gl��::�J��-5�;G���f��X�e�)���|��`��r���<���O���%�W��H���,���R���	�|��MS_h��/$">�s䲰�.eFݙ�5jOd/ó]��|���Ա/>�7��h��5���k�e"�U�� �	��ѩsZ�jiF��|b zڷ`_���.+����+�*�H�]s��?��]]�,8q;��M�,#ڌP�3�8�l��x��x?��A�j��T�]�\���0���2��ގ�3���]���G�^���7���o�%>O�y��W��,O�����l��IQ��\�n�ս���t6��0����^G4R{�*gJv�[	�9�⇢��g`�����ބ�-��D�E=��%����t�����ܼ����f�F�ͮi!�^+ݽ��m3u�2{���t(�A2�7c�y%�|ߌ&r�Bu�x�8:�ù�L�D����֤���v׏q��=��"��a�8[��msW�:����\5Q�{]�_�>er V�}�)�5toSn���@�������axP�P�����Q���*QR���P?#!���3���챭����ѷ?���qQ�}s����,���Y�|A�:5����D?�Hfǀ�Mn���0md��G�������Y����٠�m�4�-O��94�n~q"���;zg!�1�'��:ccA=`��W����4\�@����5��\�=��A����çxUX���ۮiO��������,?�������Ѣ�nfw�`a��rU�}&V�fȵ����[�aGQRE�g_�쎞����4L����O֒�-%��G�Dҧ��T������@cq��z��¢C���v�)���\ԕ����t�F�zp�����C�F�Գ�Y����o?����?�Q<�p�g� $�+vwr܁R[�����QtS��X��Te�����*�ǤӃ���������mB�G�v�UQ�oD�'5���߫5r5U[��H@�+_�0��iTxv�7��<'�s����Z%��X����t}=�S79�R��(XB�e�d�@b{̮x.�\м&CF6���K�)a�QĽ)�o5�4荊j���7-	hV�dݣT����s��*�;��$���h�=�lߨ�;�e!�c�G�u�Kmm`�2�����i�yA<lb�]<i�+�W��m���.}D�{��,k�O�P�����KU�S���Fu���u�{�h��MN3��M��k�1����E�F�$��MH������id�zV6%�<�s������^���8m��OV�{��h�\�)4-NXN��=���}��������u/�\�x�Q9�#h��J�5)�!�'�!�)ˮ�3�A4Qoz�f�sL�6����oՔB�b;�Έ#�=�Û�zLw5�>?&(4�A����t������&�"�#E�"����0�+�����j ��3�$��U���)ݠ���]ž��¬Uȕ��>�}���.��?&??���KAC2DL 2��r�qkt$���7�;	���n5�F��J���V�6��:�-���K�U|L��s`c֘6n;{��Ln�\����vK�4��r=��"���=�Q�@@���^�+@����HT�aa��[����8qkl$�1����-2�u8['�ͧ����Fը8�tH;-�
[��G��v�U}#�7�"g���̣:�>��7ne�߻�ݞ�o6 �D���`v2=��MR�g
�}}r�u�T�4�Q�ܐ����dE�d�;}!�\�@�<��c��5?��Q���.ٻﱜ7����Rq<ҳٴ�ʟ6X���T�Z������I�ln�����w�r��	+��֕M."�~P��i1&�������Ӊ&j�Y{�B�\���C$��{���kq�_���UG��!�L�Qå��e��4�+��Yfژ��?<V��H�L[�cO�D��
D_o�P)��Z�C�dʭŖ�6�tRB��2܁֘E�qv��s��_lVU��ya�ȵ��I�����SI�zڕ,~yB+G�?���7A�3�}�M�(��`��1�)�$G��.K(�x���)���6�n�,4�(�o��b����I�5�m���N� ��"<�F�S�>])i�o�t�[ׂ��P';�ڛ��׫$���b���L�zcr����D��>�;ZœP7M�Y$8����`��Q�����n=�X��6���Ou�����^�?J��;���(�7w�%}��l4˯������D�ؙ��_���5�����^�?ub�H��恷��'}7�Ԓ��P��W�_��)"^V��-�1O�	d��^Myc�ʫ'��-�f���P�M�ta��'g��\���g�J�j���Dt{� M���R����E��v��� 6O���Q���y|�Z���q�i���n]W�f�X�;�k�Ş�S8c0��h�Ƙ8Jnq� �]�f���L��q((y%E��~�������P�n�hda8ŉi@���\��V���Z;s���(q�P����h�|nX2�\�F[AT��D�M�2�W�����Q��N���!������5�@�(j�u�g)�+y�6��A�ϒ�i
³I���u�ZDU&�l��$D������Y�g[�R�A���^@�|��C/G���zH
�}~�FmH�����+/�oܺE����C��w��߸z-,�M}�S#W#=�����w2���` �Yp�H�>�������U~(�4JH�T��CV�>7>��N;�v��JZ&-W���b��di��}U��׿S���*%���Z5��6�y�TKEf�R���\�Q���~�披t���
�kK5e+���8��3��Awe��=J��Ǝ���/uJ��.�����=ݲ��C �r�ny�g���<����5��vO4�wt`T6J�ǂg�܆�TZ]�N�ܯ/Cղ�ق��m��)�,�����R��r�l�u7�L�M��z�_���Ww�n�y>qS4���-�J��y�
q�g��L#���f����X��,�f��I۸k������9m�ʉ"�W�J����q�x��&4:}Y���>�ܩ���B������3>���z��������`� D#���r�l�B���f'(���C̈��֪����u�ud�ɭ�sp>4��F�S�wH�0��5:ELq�;��]������!�Ç�[ ������
�f�!/*�O:��O��w�>kԒ&Fa�/���(��o��#����������:z��<+3S�����b5_��vds"�>��]ͷ`�Ʃ���sa��d��4˥��@��y��e}z�Ґw�N���z�F��y�rx�Q%��O&�����Z�ph�B��3&��5v�Βq����__�(:
+1N���I>Z�ҀNv�����8��A��b ��Fm��N�v ����3�[�+}��,�z�Q�?++�\���^cs�r�<a�%~l�;�E��� wr5OM�� �(�a�D��B�{��@_6���`p[5�9 �tK��-9�ԚJ	(I~� [b���4fN�m>����^����9�9���]?�Di�*���a2I[G�����m,=���	�t��9����7y�k�,^ӓ�K�.���i�&q�^yxj&]E�u��+>r����7��'uR ���+�c�}�/��
���eW�?"l�c<7'�7ߊ.(ڈ���+B[��vOcP#��,��k��R�,e�(��УU�L�ۖr&��(Uk	C+~���E�{�ad-��Ks�������������e^�ioi� ��Ro���G�ѕ�,̕Z��P��n]�=�oeq�Xm��mJ��j�ՄN��v�/>νa/ΰȫ�|�ᧀ0��M�V6�6{���t�("l��q��(������M{o�l���2���>+#K!���8���d�v-�kp����실�/饸N�"5�ՖZo��N�i�J�\���!��פߐ��=�QG�K >�VHR:�@T����(�#sy��䴥��������� --b�����tV��4���_�ϱ�nC��9�9���͍�Ld!o�@&��&�<��Jl��3]��)�3띝��{9�M݂��j'7?�;�\@c�� �|)�������vk�|��%U�'�{�weU1��nI���`By�a�N>�}H�[i�F�i�cʊ�Qr�!=Lxq�Y���Q�	�6�k�>ASt��#�Vx�[�_����rM���1�#�j�D�����$}�&�^zhCH�8G���$ߙp�u��2�鱘�	8�w��5��n��K藪{��5�U���,�y�M�ϫ�ԏH�l1�%n��W3o�G���T���S@�w�9���L���^���p���\ݜ?̎�RWk�lR�v&�1�f��J����t������"7R�}����~�[_ZPx���0��q:'��N�H�ƴ�޾�0����6��=]b��oʼ��T��3LŇ�y� 27���$��B����Df��Y<,�����8���+��,j�qF�DltA@@@DzSQ��ti�.�@Bh��#M�RH�D:(�БZh��-t�'�*~�����ȳ�^�^k���k�XSˍ�8�˚���>>�4�sD�������jp�d�����~��g1���Q�E�''յQږ����1tr�	����tw�P���%['�2=��������������E�:��܃�����%֌Xk���<Op�W� M�K�O��*ś�@nx�#P�G���P�tm�^Ng�0_AJ��#m���c^�zWH0`%��@�%y$�iלP��#`&��h�,CGQ���b�'�9#:��|g����6n%�l�in���ww\&�0K�I1K>Ϡ��3D�eM�������l��_�:b/?+]Rz�^R"�mḩ̌l5���A#˯ uzX�m���C��L��0@z8䬿���J���S��M�Ge�N��G�\�T�EV� !ex���e�#��P/Jf��� J��,<v�����D棤W�?&�'VT��p�hnG�kly�d�"��ɝ��Tk����d��)cQv�	+�!������r�C(M	A�+�r���O�3Y/\Т��a����� ����8�^����ߒ|�Ȼ��sHR�����b[;b��m<NȦc<�WNɾ)���)<��&.�Ȟ����p��� z~n���=���x2J2�@���	^�Q<���١+��T�]��j�q�b�6˫�`\e\������+��}%~����=�<�pƖԑ�P3��B�?����pw���ւ����[����~t�R$g�g�զW�db�⩕�CV;uu��?aQ�d�{�eb�3�5�@@|v�d�҇�y��[%3�o#�N�����#Ȳ�;ճ�?nٚhW�� �2�#v-݉�苛��c@�A�V-^�b)>�;hm�	�U�Q�c՟�B���ik!߱��v��X߫�ͼ�ŷ�8�b=erY��,=�xV�ԣ�p��z�־<���/t/V +۠Q��?������Š���"�\�������=����c^:ۙ1&��l*1휧�	+"��W)��p�c��Z`]��`�dfis��O�q���7��ٌ��|͓6<����ՔJ�����zY��t$�m�?��Y��i���2����#-����\�^ͬ@=���
��� ̞/�5��A��۟-@�tAO{`����(m���K���gS�A՟�F	�����t����Uo��Ip���{5���	� ��,`E�oTֿ����0 F{�L	j���-���BGs'�\��Y���n�_�,�m��㇁�ř�2d�q�M��.�Z�O�jrt����R�US�� ��~��Pzɥ���.D�*�6�+�u�u�F�>��~�ɓ}k��j��Z^�rrPׅ��V7��}��J��h��k!qXd�)s.�%�(�]�늠��,�kg�ɓ�P��t�}B������2�H�*���2$�񈿜plN��\�k�#k�ZD���6:+y��+0��ТЎ^���� 3Xm��6�U�7q��dH`���D��y�徵�_�.��4��(3��:���	�dU:�����g�t�P����i�v>A��2� �(����/�z>�6n�e���!e�����pg�"��ͽ٢@d>��|���˚�L@���A�ϐY%a\�����΃*
�������V�1R���[�҆jn��e��&���i?uwq���W�ϠZ�`:Y�p����z��2���p���l�ԍ̉{�̕��ͳ�#�z�!Ry�{��tc<�:�X���w>C��x��E#��[p�#�#�|u�����~^�����t^���H��,-���څ�;	��֓�e:�h��������0&�/��m�@LY.�K����?�i<�����Aqz�lOy��U�S��l�]�ۑ��%���čg��r�3d�7��}z�NG��Ǎ���F0'p��y��ѻE2����� �]���{�з7�%���\�>�I��v��/o >%<�Taƾ�y�f�)�9��/(���-��kf*�y$_� vI ���(Y~�q-�n���&ɡ��(���jV�?�|�r�kk.x��,�<�oZ�%i�f'�@g�~}q��!�#�GK�:/�H�o�M�o�+�"K��J������C*� ��G�Ј���lkZ�'I]����;�,^�w�hse��E��9gي�G5�����4��x��u�� V�B�z(D5�44k:�Iv� ��ҒX�|��s}�������'�б��7p���ҹ���2�?H0S���x�_�t�a�i��������Ӓ�q���W���~<�$i\C��bh�ju��_H#P�a�ܖ�G1ނ���m��D�3������qW/����/��G��)���ck�*Q�&'��dG�[Iۇ%����N���k����c��g��r�����#w��o6:$�\�h�,!
���2�o�%�ɻ�w��Z�cO,7��b�g(V| i��Ts�ȋʽ4z���ѬUv�jt��'H1�Qk*O)��<�{��|֭�u��ENI�5����f�G-��շ���v�a��Ǵ�u�C�\���;vߟr�+���$��׊5�=��j�����u�@{��.����L���s���	�Ny�B>�����טYF�+�]\TR��� W���\$ae�3L.��"��4�E�#W?<ɞ�Jl4l]�hI4�˝jU7��>[H-Dڢ��;n�|w����:����#n+F��l�D����r�Į�S�؋�h',:8�K�	k����d�J �������髿G�u��T�F�>Kz��ϫ'�/��ˏ���+�;]����|M��x`)[Q[K�~䪦�E!f]
$��SN����E�)G����A��r��ړ	fA��9憉Ձ����B:���kH�ǽ@�C���
� �Zj,f��a�UO_����c|®9�v�h�c����ev�]{���׆1��;�5�u8]3�,�f��y�ێ�K.�oiLI���?����Ox���� �ol����^q��9}�-��|��p�,I����/��K�gQr_�p�1�|���>��|K�iӻ�/�Gފ�l;���Ħ]L&���Zk\'e��ݨ�~bVuGdu+���V��o�*�{�!��M}_ R���n�%!=�U��3@m�2A���e����U�י��j�XW�N�Jl�-9][��K�q�B���,�*���J�K�A���rĽ�H�9���E����I�^鿫�̋N��$LNM
Oy��W������~����oFW��Y� ��o�	�v�5K�Oڊ����Uڌ���u+�/;9v�n�)ޗDw�6���]Rx�<�?�M��}J3��#�I�yOn�_�1ę��>pف�Ұ���<�uϤ�nL>Q̈�ڟXͩ�5�^�s��qQ�M^�qY%�/{�BT]�7W�l̓�)��P��H�����7��y7����O��;t�RixB�j|��K�2V����ń�̣$�.XX��0~��٨ƛn������ﰪW�Kw(i�n�B!�����)u;��^:�n��ą�J�k(�sˉ�)����n�'�e�� ^�ǯ����ڒ�`Y�Ij�Ms�Aō�.�kĴϙz��6s�͵�������<���H�V[*P�z%��L�(�v�V���R�\c�93w�D����u���p'9V5��ۚ��FF0&���dZBgJ�9W�^��b⩄W�ho�ET�"r�QY�':�5�5���4'�S����u �3c)~� ��3�-�eq�8�g���СJ�����6O�Z�FZ|��T�o� �y���� ���#yJ XS$Ie\^Е����� {O�c��J�Ҕ��g ;;�Rӣ56�t�~�fS�+_�+Y[IpsC�k���Ý�u�c��,C%�<|~�J��7����Pu�4�u���/��	<��/��K�6����~gm���/JLw�׾nl�GD������3�#��Rw�Kn<�>���u�D��"��t��{(�*tcZ�D�qQ8~�s��\�Da�S�;*n����ݤK�L���۝њE�Gݴ_�Ƅ�^��~�ǋ�b��4Y����N2ɒ��Ρ5;��n��T
V=5h�e�����,�y��HF��}��}U���@���h�#]�oƶ���VMUEŶ�����yw���������iE�������ʏNH��q�TnM8%���>��z��f|���B�
���?|�F�׆���j#��u�wn El!q"�ϴ|
��{ո0v��{]В�A��H`����fO���{����STP�[��w�-�[�a�Y'���X����6�,�T<4{Y:����o)���>]@ �;O���ۯ`��p�}��X�w�}�Bh�D�|u]Y\;�{��R��']o}z2<���`L�,�粈j4G��^�A 	6ddR=�3�4��u�yb�`qAN���m��]�i�:�N? J9����H�F!�y#	��[��F E(��	�j[���S�����(���y9���<�4z�j{J���;W���s"�ƒ�c� �
��ɚ�}Y� �n���~η��f��k�8�s<�&����?��Ҹ�����Ilg��5nñ���Ľ����g-fW�V@H�Ϋ�/�W����ٛ{,���ZR��{������nvL�e��uwmDU������~�S@��X� �X��zRl�v��9��ݙ,��q�Y��Y�E��4%��ps �s.,�@96L�Y���=~��\���8�� �g�8!�]H�SD�%�4���|S��E�);wїz�]b��;�6H���#fꛦA�V|A6df�~1�����v�V�����C��!&���c����"oZ ��a�E\Ɨ����jS� �G�w�tekq�����m��<죾���e���ۇ�/:�7=��(�<=7�|�p��	�]�9�������'nAGL���[�3�wrތ˲��5�_ѢxD�?n>�/��d�]4@��4��v�/X���%����w�t��!�o��*gL&���a������B�G!8�8a����-�z{��(���˧r��QlJ,�����P��������Nnej0��s�����a�- �-w$�����NE��x�HKI�Q �����Yĥ �D=�N�<ٷU���1x_k�3�ë���
�u򄌹�ྞ@�|O��v����ˑOp|9s�q�O�Kq�<i�h����7y�k"R�@<̋DK���)>`�v{��Y&��#�x-�wR�?�a͋hd��ow�w��.�s2�����<�n?cb��0��b.�t�X럠��}�9���4�*���|͙��f^���/�1��C�`�ke�gwjzc>9~uu�"i�y���>�����l�G�LBȢ\���s
�ԺjKR��`�x]��IխǓt��g(�R�o�= v`�N�� ��m ��P�@�5�������7�;�FD*�V���++�(�q����@T���u�(�(��h&����Q@D�	�Gʙ.n~>2
Y��v��{�UΘ��X��Mt�cM�[Uidq�	��b�Ź�4��yo/����S:e�����z�}%l7�y�z�}�>�.;���2�:���Mʿ���wZ�d_rn���aiڅ=ܾ�qvחB�N{ۗ�y�MOϦ<���H{��C�����y7KC-��d�.w�)�|����-�^��,��������֌�����D�~���@��v�N?�Ԓ�fV����oS�uw~�_����ѡy�/���
~��}�#Ӈ4�d!�tHȓÔ�s/1��G9w�(�e�SG�u'�Mqv��>�feqc��1-|����v�J:<U�*������2��+�h��<�u"�: ����k�إ$48&��	)��\�
ٕ����͞����Q�V���{���������/�s��oC�>$�n�.}�-k��D�oJ�:��ɟ���;kJ2NGqs���V�&��r
��"���B?N����@w�ኦSt�|��aY�Xܺ�JmN}/Ͻ�S���䫙�:�R��Q�z|l1Z�+e��j�;̈~)9��?�#ETz��!TY�
�ހS�j�O �xmE{>V>uFY��n;�L�qnݶ6��]3ܗ1�|��g���4�G�|d\Z�X&�W��%%�dy�ֿx���E������|)���ғ�v)(n�X��Jf����O��M�ۧu�&�;�������w�����H�b��xBNש#ؾ������1�B��j��c;���4�9')�l�T�ň2��ӡHIz��oE(����G�N^�(d(�_��n1�T0o`�_2帰�F�Q��qQ�x<���g9%�6|�U�Ã1( �s��>�%���U|�O�g��]č%.D�Y�Cr)�ɕ�z�`�er���<�5����Msh�79`<��_�л_]�Ȝf�����OM�$���s~o��0� ���{�h�T� �RT��.��
���%^���K9�٦�K�{�{��-�P��r�C'5@3�dOt�ª.u ��%�8����Fֿ��w�|�y.�q��U���G��^T2���<�J���J\�p0\P]*��yKV�-6f\�d�6��0���X`�?�?�P�H�O���	vЈ��_��N�VH�\)�!��8o�rx�O�R�߮�|gہ�rI	�p��՝Oj�Kc������4����^��c�~>A�G_��P��\��A2��>��0P�]���T��>l���+E��Kڦe����6��;��]�'��ȬvO�f����ɹ���y~&O|�g�em(]���"� {���ʺk������*U�am;o�R�?�9���WpW	O����q��n���o�ú��x����s�����KƟ�.���P��(�j���L��^��;�����ގ���s#׺齺Jo:����؆�G1��Cߔ�VD�{��x�l�`�ȳ(��H���W9ӳ��B�1�ծ��
\}�Z������ C�������#�$#_ހ�E��l43�5�Ɛ���L�5�æ׉�U�,�޷� ֒W� j�t+������ p�G��t+�4��ȡ���2�$X��k�Ύ���1�l��ɸ<��� �Ɛb����y{�G�߼���׶*}�چ#�_��P��}���R$'f8*��+���!�R���8�<��x�����yO���l���݆O��fm.�)B��$)C����>���Ջ#���{>Jv1`�xUee��' v������!����	>����W{ޒ��ZQ�����ݻ_����ߗ��h)e��2�!�a������^�h��f�B����W���?Y�#�1&5eX��>/1~Eܚ���Cj��^v��NDke[�bz�j/{h�l2����]��nu=�C��m41�)B��TQD>-�݇w���� IM��ߴ���
H'����L�߅�5us����^G6<!Hi~����m��f5����H��2L���\�1�-�a��gnƅI�����5G7W2L*po��W��ɛ��4�����c�V}Ȳ�
o���-H��"5����R6�0&�;C7� ��{�l���w��B²[��d�$���Jڟ�Z�z��k"�����3{-�~����N[�T��qR�74#�]�;�
5��e��{sj���9^e#B�x�e�]4��*�B�V-����}N��fTx���:E��1�'+9��⌁���¼v-����v(�N��Wx���@`7�MfY��]2K�v�1���^�te���Z9CDDv��cV�n�[������@���7#[�9�2�:OU�42��{�-���c*$EY��A��y���c�^��~^>��������Y�1�2	K������1/ٲ�S����2����;떗�}�I̚�n�ѽ6 �hV��Ҿ]e��q�y��̗Q��9�(|9#�#l,,r�WK�I���;|��e��"�����j
,��| �oTba3�u��KҞ�ظ=5B;�T�� �5�>�#��j��Q�N̠�nEM�ʻ����h�)g�
��o�dV��+�(*bI��W���^� c�͏��$$�+]������ˮ�~�C�u
�F)����E6�'I�z��S�6*^Bx�bl����V���c�FW�2�!���ۙ�2�n���M��v����_�v����G��䭄�jv>]�K3��;��l)2�7���e+���
������p뇶l��w�M�{=�o�N=.iF�Ԉe;Q�v*E��*��ᓗ O�#�4�,�U��2u~�|];[lF��b��!�9~�oV��%x~ebo�Bq����6I'���&1Yp+�F�W��lc��c\r`w��| <m
"�o:Jk�X<TP6>�����s�;�W�,w�������}��������kP����ԛI]M�4��Z�O}����A�8���澥d���`2W��Ȯ�^jŀm����3[$�	�t ��v���/�6Ñ��:vɻ���{d��ҏ�^�-$t%JED"TQ�-�g?8�9��"{t@��Mh��,�ڮ�ݚ�6R����5�����9�TZ4�\���p�e�2����N2�w�<�4�o��7�;�b�.��*σ�c�	�����~���ÀC����l�Ҋ��#�2�A�l��X���d���J%��k�痏�>�A��={��ۛ+:Q0�����>[	\iY�2�5g(���cS�� R�0�x1��t�-��栕%��	�	�{�BJ�`F��y��b�����|�^Nɻ�a���!���i�7��7�$#��K�����MQ]{�;�^�H�G�)��D�������	�����C^��	�p�{��N .�5i��#"v�Yt�
k���L����.v�U���w��{��Fj��� ��(6��M0�X�W#��hWg��Q�H3.�5x�Z��W�V�ri��/�<t��/<���>�ɚ	��0ٳ�7����BE�L�I�N(�ǘV���HꞳ�R�ܤ�z\iD�]"�W�1mPdn-�W��m��?�NF%p^9&�mX����R�I�t� ��:�hJ�VԘ�'ܩ�Kg"��Z}xv�ɴ�eC��;u ��,�y�s��"׵>�b�s} �9�������`|臯��3�]D��#��rȸ���T���}�hEfs��4�ǖ���{�j��kB�L�Y4�'�?\?�X��UW�a/�7�ks��2T�ݯw�ӂ�m��cK���8��$�ܝ��O�$
?��|�j~�#�/h^�����2 �@�*����_����YMw�׍��K8{*p��\�����`�����@��������c����^��E�^��b'^"�S!�0(9�Us1���� ��I�krk��z���-^��k�᛽�1�ad*���:\���� �q�ܹ����}G�}�+�/�i������Odk1�	4w�����Wi"X|�ݵj�x�yh�F�|ߨW�|fh#
_��_R�gd��MnaVhY'����#f��J��}4�x��TD�&�^۬��@)y�Zs���t�xw�x��n�#M�����:�d��4>�����]�x�>�7֒��)��J�B���}o�h�V�X!k+�/���CT끡��K֡�K-;���nx;��1����|˽�c�ɜ�P���X��JY���J�&HJ"G����jоu������W=�����h�]d�{���֤Ny=���F������2�X��&��]I�t��8U�J/�^fm};���(lzS�E)Tܺ�8��U��DO�H�*�c�{��l�PF�C���Q�I�MY�s�lV�%�L E��(ĕ>�f�6�8�jｊ��A�������̆H������bH��p�˓pM�̧�X�¶�s��|%�|�Ȝusc��@]a�#���w�RE�嶽i�|�1e��eA���d��NrĄb4D�$�8��Yl4�qd��^n��0���Z�j4փr���so����^����^�	���}L�>�+�,&��Z#ӑ�o�/g�!J:GP2�V��C��l�ƕMYs/_�%'�X%��EV �Hd|���UR8�	�=}�\!�!y�M��أ��n�N��/nƧ���.�(ź�r�h�]L�xSSP�h]�(f *2聽���@�p;�w���ķ�&�Z�C�m^�\��D��Ț��/��J����OOrw-P���e�!���M�Y��"sr�>";ԥ:�ϐ_'fG��N�[�rY����\���e^*�����i�nn*&C�.E֬U��ͫ�Vt^���Y�:Vbߍ��J�(+�[�!�?C��뺏�H�E4�eW;ʖsŅ�7��v�,^}w.E�����W��h.�u���5��Vr����}Q�A���212���̙�M#s�&�q���d�:��f�W��S�l���`�ė��sk��#|��麋�1'MT(xش�_���A�廲�F�f����>O�^�W_����o������N�Ds(Ją�">Ď�[tT��e���'���u/	��OӐ��h�^�,���n_��lޫ}���4��e}ޝ��V�$&z�c�S�K�-6��bv!l��p:�^�ǹ�2�~�j|��^M�ػ��}��D�8���v]�\�E謊a&�1l�ˬ��4��~�?�k��|���Y#"wi�I���/˖� 2���Gѕe�R?�Yx�D��K��2��(%EsB����f��]�ǫ�"_��R�����:7we)r��ً��vB���׮Wc ��h�[v;��e��oS%�N���R�Aη����8:��r���j�m���=���,N	��ފ<��47
�hʼ>��"����T��&�p�,�f��y������De��\gu�K/YIn��׽_�E�� @w$O�^QW���2�@��1F3�􃓟fd�ܹ�P�
�hٟ��v�������+%�Q΢���d�;�x-��t�w�TrE�[A���N���F��E�`{_ҹ�_&���$(�n�n~�XL܄xȍ���w�M�n-}Ѫ^؉��[��U�=�����_���J�l @}���b#� s��k�7�����x��Ce�w껇˦v=wH������E�cϪ;���������]owP�W�,5W��|t��i��#8iT.s9�}�{x�u�&�v���l���}��7��GPV�zc������p$�5��[����vF���[ʆ�gj2u���U���-.,I��x�����c��|��br!�ËoY!5v�c��p�w6h��r�Z���49K���:���p�w Svy��-���2��� �{���"|�zRa��*����G��&rl���S����d4��.�>dd�H�"��)�C��H_	�l)]���ś�1%�VHl�7��&��j�|��k�^��>O����ɇ#�.�Q�;d�H���[]������XvL���xjc�H2���K��.K���*���Eσ���=����U���d���v3f�I�}V^���׹"�,�y���a��o�0����u��[��L��%qG���wj_y'� mc�޿DrX���m���,��2��Nn@�	Q�p�R�_E92*���.{53j"�ۓ���d�lʗ
^Vz<��R�<3�/����!�]���:��ľ!b��D)k��P��nw5�4,�#d���
�����g.YU=���vu:��0�	u J���� me�:�ZI���+a	�F���\���ߵf�����Y/��f�5��D��Z�'��ӥ��o�DJ����^�YeM�攗%>{��<fN�'gTV��1\El}�$i626��^uԪ(힔�$XDNn�#}����I���
�_f�ɽ��b�C�A�&�h��[�;F�r�����f�t��B�wj�M����	(�M�!�dYT��dZ$=!���ӻ�C65T���֥�0���}���lb�|�_��;K�r�Q땦�s��� ��o�1`�j����ڌ��2|�ܞb��K$����aG��ꊳYn��R_�)zm1��b�Z�����d*D���t�>�������Ϻɍ����#IN5G����2��5".5�0�./b����D%�vX�N(76���U�7-��뺲Gϭ��y���{$I�:��������V�ƍzF�9vǳ����9c� Z���NYrb)��'�¶%����w��/c�ݠ���G�%CM%o N�;"���GH�[C���A<Z܌��|M�����2����S���Tr�������7��sQIѐ��\=K%W��Z����K߰�@]+6�o.2�']h�%9w]ZJ��4���&6�X�%ڧ�V�/������2��@�]VF���k3+������˨�PA�ʛ\"�U��
�]��nfE�y�i�uC��l��뤫��]�����e7�&��r��[痲��>�y���D�K���NX_�&Ķ���v&�׆J�s�hxw��]\CI{�|gq�� �������V��i�b�_�bܪ�_�;A���4���J�r~�>��mW���c;.�.N����c��0���+�Q�z�_��U�P@>�j'� �ti4�r���e�p�R$��=���m��'��8"�w(���|�}����ʣ��G�o%��7�$4?�?���S��U�iV���MQq�'24��y�s:[æ�\��d�1�c-�T^~�N�k�	 "��g���}F���~ۅF�'�sױ��s$d�sy����̗��٢7���� �k����6�.j�ܓ+�H�)C�	D;x��4���p��"[�x��W�5�;���Q��T�;h;�~R놕�&$%�=+�23���N��]���\��.F�胚VĉD��v�A2����%5��ؚ�'� \��v�\�����F���S���<l����Hݍ_��d")@�Mę��`�T���Oڸ����{++�i���NFW�5��r��
�*�&$\Ue��k8w��%��)cW>@d<r��I�l%}��M��Z�R�8�a��
q)B�@�r�:I�����J}s|�`F����EXa��[�Ee	�'2<�.)�5������	V=�<��3�W�
	!o�>I�`�J皋tm��cl1�1v��Rc_�4�)\+4�Uhz)
��%��[���(�ATd���MF��I`l݊A���*>���d�b����Ӏ��`��(�.����P��U9���@m��)˟�|���S�V����@��{a�K���e XC���Y�x�ڨ���.���{��L?���3�z.d�)`� g����ZI�P���G��`� �-k��K9��WJ!&��L��yb,�ᅬW#2�^�:�J��LW��1*8&0GÒ�ͦS"A��f�=x�WD��*==[���{/��T(Q���wˏ�����K��ԡ���@�����:U��r?�����@�J�<�0��h{gnd��j삒���u���������xۉ�v��ɭ������O�1N�tC*����Q��������y>DP8IU�����pO"�@ї4�g�Vy{Z���8�'A��D@�Ce�^�S�	���}ή�H$t��-�GE����?���W�'/��Kbm�╩+7?hx�hU%N�V�)���#`���:�;^}��B��ϧ:�+���[ؘ��C��KXb5dNMvS'>�2������q����J�����{F'7���QK{�M.��Y��1"�>�e��s�h�\�����_�A��ӧ�kd���Y*,�Ҧ�ɌN��_V�j��?��>��y��2o'*�41>o�_\�@<c�wU����ڔ�߾/R����ԕ�l7	`(��	͗,����%Ēu�ߺ����|�t�+Z���d؄J&���ΫIl���*f�}`�+���̬xç��<.��L�(�\�����F�F/���w��˄��2�a���fe�|�)����Sj7�y\���`e���Y@�N�����/iΚ�2��6�$�bΊ�*2�C7L���y@7��,��p۰� ��@P;��I�o	ղ;a*�` �..��<�0&|�e�-Fk�$z����R\�a.��U�?&Ӡ]���*�����G�c��U�N7� �/�:6R"
T匈Y�^����W����>�N��*�I{�ʇ���в��� y�"k'%k�8�R�����6,�MR�5�g��i	��j	��7NU�<�Y �����5�U�Z��=�ֹ��/A�`ݾ=)�&O�ơ'����u@��0���SA��<$��K���8���� ��1��ML�_��#+j}jz(c�"�@�+��ǯ���%)��k�PA���7�S��[1��t=�E�:P�_~��T���:3�QjIŌ��D02�)�Q#�3j��ٚ¥��|���A�E:�9���N*;=���>$������ �u!��*�?&��h��M�dA��st�=QpKX��h�7@K���M��`��,���x�ύ\J�j��J��Q	 g���y/�r�n1à4G ��4(�J�!�:F*�$�^�g��cVė�eۛ-?e�J����\	�<����������+��1�JIe�j�σ~�rIn�$��K�J�PKv�Aq��VD�c��u"����W�1�G�����5!�nWx֖6#F~410A J3�7x�R&�HFG4�(��b���w��}��[̈�f�t)��g��(G��s$y�Dw�� Ee���(;�QB6C��VL�~�[�رf	\���Ɂ��b �H��8��o�"����&�ߤ���*72~)����Ç
�Hb��z�1�ʡ�b&�wJ�S"0�?�V��i����XM����\aN�+���+w�V��J�݃��8#_�͊��V��_��	b�/:��bB�6�s�1�<c(��O�!p�HPm1�w��oZ���"7i..�م���}z��ݣ{�����i\�c�"��|�=vhj:�z���al��¼#���yF^��o��|;��1�h��'��=��Z�'���|��ۄ�XFJ�+g,��@�P������PX�+��T���b��mݖe�m�w�F���jWÂRZ����W�"���SϞ��/��w��ߜĳ����#-,�������l��������_Ϸw���|�_��O��� �_N����K���_�}�9����?���} A����Ƶ.Ϭu�)氺+���z�ؽ�\���\�����K��C������T��n�ogg�́��[���hRy�m�$O��A�Z:��W�_�FRfT���"�c�'0� ��G
���(e뱉���7�G;�%y.|@��w{A݋S��T�["ؐ�گY��h�:,��:�H3��OىB�?�,��0���>��˝5����?�� ��r̀z�62�a�%=U;�W��
HL\i@u モ��52������)��������Z�/�ٱ��̋�b��5�+-6G�
5�����mUv�iU�j���������ӷ~X�y � �8���+̮�R��6��buu�#�w'2�����,Q�_u+2Kʹ)�������e���-���mDҥU�2y�Ld�0!���V	Q��c���A2Q�N��֠�6X5]�Jx�M���3i� �{��F����}v�aoq�BVSp����BHe��`r�����	/��ێoJ��U: ��;:R�u��������u�eyx�a�0�+R�T'z��S��ɧ@����9>`>��(_Q��a��Q>/vſ�N;�R�7cT�^�����1�s�)\�� Ȥ]��W�t7w���@�h��B��q�VG���Q����ny@-�g�����)Z�U������	7¶b�j����7�W5ͩȠ�����������P&.��=��V�M�]��Udh�y&N���w�?N6
�� ��.Cm�H���� ����f��3�I:8��������T�)���.pN};_�#�'�hM�Y�&��[;��潌����P��4]W2�D�:�R�������I���X��Oo�(J���y�륂>��K�����!vI�jyfgק�m�g�/�N[��� *\�/��ч��nY��� ��*�v�*��D�%�=E�^l�x�qB�p�%KL%��_|VW���(9Ww��:�G�РO��g��3�T�'���3�RHj����'�\�
�nZQ�N��]R;C��/��Q�+|/i�q�|Iw
ņA���������.vVsrp���X *S^V���������X��
�8O}OL�=��]M	s�D	��M���C�#c�뻀z�L�!�m?��9�)�n�{���ي���0d���^��m�����M�jxB�y,�nH:6VJ���]r��&»��k^���6Q���b �O����Q�\�sq\��P��Y����Z-B��v��P�d/���V..���fwJ���Q��G��ռ�X�(�_�#iQ׶e����7E���k$~���!$f��h�d�x��>���F:� �l7	�Y�0�6��Y771�0\�Lmq��������7��i^���:�슢+�x��s>f2@�z���r���3�*Nl���t]�VǶJO3WQ�(�7^�Y.b#C��^�ȕ�52��ɒ`�M�W�4^?AU�iw>�(\��q�ҡ=HjZp5�|Ѿw��2����w5�h��\��|�p�ms�f ȝ�D$�l�D�������)H��CpW���~\i�9ŗm]Į�5�����a�N�#�ty��?����v�h��=�d�����+Л
|%����~��~m���\��W��N��O���Α|}H�����
��f�z������Q�Φ��GTn� �� �J ��Oz(��@I-NLp:&I�:LB ��H��E�7M���IL�����W�3YG�~���#~�f�~�^�,��}�c A�����}���E�$6�'�D4��1x5m�726iu=�}s��DA	h����C1c��ws^/g�:��@��W<�����G�n��鏔Ñ����A��\�oR�*� J[K�v8d��K]��V���+٦~OkgLd�ifXh:��]W�D��bOK���P���a���=M��cf<�\���L�>�����
0�?b�ii���a�WBs{6I��/G�z���)hE��p�&�P����VE�}{ۅH�ײF1�dɾ�������Zv�Q�mP�gƾ3!�����|��?�t'����k���u߯{7t��@�smT��s�Ǿ�7ý��z��Q�xz�7C�C�Ǚ�*�9��j���Ů�t�����k��������XIK���쫍�"���*�\۞-s]����N+��#E��}R�}��^!�4A��~��2�	��K��"��MZ����gFRN�o�j}2��&_?�Bja���E5�G6�驶�Ȃ(� ,b�gB�FA��/돓Hn��`�넷p�-~�O�$�&���K4��#�K�B��2r���LЀ����?I�\�V�#ɵFw0�lS}'P=�.#�����p;��Ј0�"��h�����b��3�)�Y#�Tw~�Q#�� �x�}��-��"gF�
����{�^�Iq]��(Vi���O���4�b\d3I�h�/���ۓ��O�;�# O#珄�V�o�.е����J;F+�3AKE���u0B9��,��URRY�A��/��t[q�a,p9�H��啕�U7s>�<S�����G�����4�}j}���$�a^�ȏ��4+O�Vt-V��*�x�',�%	����J�hNr�5����\pnL����5G1�3x�'�Pl�O'.���-�ϜG� ����wR��PR����5'Sӝ]1�܇'.ԏ�i�XR8ACM(#�H�)���Ǉ�	���*�(����?qW̟z�<m0�"�i������p?|X'�;�3�[�'%ʝ�Ӻ�}�s��b��H?�ւ�E�ԙϪ	[��0M�nH�O �h棒�ְn,< 'R�vC��d��q�J���	���-��c��vK�o>�@�{����VL��L]����z�����ia�<���/�J�c)8�=��1"�ѫ��c��1�F�߭�}�[�������p-�6�������!�H�i�W�am����h�����yJ��E��do��í����V���+1]��=����]E���'��um�;κ���ɱ!pK���U��0�z΀�X�\��PՔ�T���i4�7�ۗ��2ϥ�Ҝ�����p$�35�@��,��e���r�Y�Q��Ћ4�a�a�5����0��LU՚ͷJO\��L��3e�%�^�>�׀���;p�@�"�H�����Ko�l��	H!mjE����v���DT�c:|T�*4���I[/���g���`.@�?��MHmX��x8Q�6�9�hk�"�=�����e3dW�0.��|/Y��w^�PѣzCI.ح��짐!x!n�ЏV43Ӫ���1N2nw��۳�]�7�)��G�35.L-��'FN�("��s���M�-��V����5#뫜��-ǲ�;�u�7�a�5Bj.�#��R�cbzn9&q�Ep��}(��D�`�nw�6���e�1� n��������L�?��T�Q�ԯus���昖��4��đYE؟5�b�����6ұ����.�ẾA8�Uᐚp$��n��H�ظ���O������YR�b���s�dDƻ6�(/~
n^�)���RAp����U���Sdd#O���� �e�:s�$��c�f���U�j�Q1�����F�&���vզ�|���D�3���u#��vzNQ�-�ٍu��=��6���7Z��c-��dk�)���f�?���b�Q�&[���-١� � H�7�֒��(����u�s�@�g�k�wĎ�M��~9�暴z�76���&ǚ�襆�);���
>,�����s-ĮdF� ��I�U����b>W�М=���J�c��m�XZ�_��M�J�ʩ��M��;�"��3�m�OT)��E�K����?�wYJj6!����I���a�Q��G�
ԈteW����0��W�WT�5�������A��E�"�*1��T�T���A0������t����xݒ�ӞՄ�3Xa;�8H[��nZW�؈;d��D��:6w�;��ݳ)�ӛ�&�+�P��1�a-}l�drӆ߹X�2��1�"��彡���k�w�a����H�;N�H�J9�t�����T���!yF	�)��Ԧ�Nx���zm�g3�6��o��Lu�(����m0��7~�DL�l�P9$p</�۩��Y���l:0e���8��R+��t2r�q1�A��`�������k���\��f���v�;S���
�2���@��eR��-�4J��KCE�G�W�r�8�V)}����p�lCs�h��>����F�*��	luh'�x�`'�W�v!y��۷���L�U�@`�d�����*B�i6��O V�b<��F�?�-�>M�눌�9�b�	�2�,�tD�E.�Q�z�f��c]�{kkt���[�=.܄��8�o��������k����np�_�s�N�I���o�]i!��|�H΍&�H}�J�3&�s�� �ܟVa��#O��U�3�#=)������6w�+b�"�!C�բz�R��:���)z�����k޼\�l�M��ֿ_��eN���&|���l���?�"O��EeL�&mb��!G3˾�G���:'r�������r���y%�
�uw)���+/����b�ޚ�`���ղ����s��b��jD���je=�»��"1�����	+m�.���yQߨ��\�t0x6.]�����/����
�μL�t�s0��S��Ö%+EԜ(�?����ձ�k:�;��v`��mg�x.���������"2�!���'��0�~��g�!e{� �l����m\Fqs���X�>Y/+0��t�ct<���� ���N���[����
��3E^�]]9KmW��a���N�r[�5!M�O���z�Tbnkұ�N������[6�=�NFf�U�{J�v���"��Et��z�рl�[õN�Y���U���N̚���C��q�k6��<�}��2�=f�.�۲0?eL�]�@��i܇5*ح�&?����Q��6�tWLd�V��Z��z���>��"����6��E��:��bV)�D��h$;Q��\$�Q%ρ���I�j��Ww��M�y�%rwV�W����F�x4��k�,�M�t������=
��l�����?�~�>�8\Z�O?��#H���ݠ���@�K`c�[t�
���4-�ǎ���KWK��
�uA�¶��]��¯9z�y䐗Q�>EESo�70%�8X�T�[6١
8bG�r������ig{�����>K#���3v��)D5�c� )R!��յ*��Y��KJ��{G=T�V{�9� ֫Jd���u�̧�+-��;�N�p:Ƴ�5���/�{��/h�ↅqCV��X{l�k�"@�"����ƱEb�UU ��\���-H�cq��2��\���*C���>���F2DP<�,w㏕5ew�qc���T��j��f� ��mG����Wa�1P�Dİe�2��h-t�
D?醉�GL��]J���~��ҶC���>�H�[��G5h���8t�|q��o�m��tu�%T��f�f՟j��PHzٟ���mZ����h�^���O%t��\M�6�zGD9�{2�����ɧ�_o����^�~��"-�: N��?(��4���$��Z���u�6 �A�bxW�r�P��<$�b,W��A x�aG�V�`�������Ůڏkq����(0�v�E̍�н�p��e]��ďGV������\<X"�V|�! ���}���
d�ս-�Ñ�� �[�Q�`
��nbU!B��	IͿɓr)�V�5�2l	��?ަq��|>���zb��������p�Q;���5#�Y��ǹW�������Î���3ck��>��
z��ހ'k�S�j�yy�znk���M����lu�)P�&S^ZJ���[*>~2>/�QaRՒx�yC��o��h��^����`�[Y�XU��ts������!�hL�l	����@%)M��˯J��h^���w!���6��J��'�ax\P+��@wk�\[�=Y�?~�%*�|�̞�Ș0��2*�۪x���Y�N2a���Y�d#�#�~*	�>�6N�}f�o�@��9���k�M@�k�Yάel������k��4���U�]�M��3�\���ǂV9���̑�zSZkl
qfo�jU�e���,�/�B?$
�߸��C_v��KD���D��S���(�ù@mߝS}-�ma ���ho	DZ���>���0�Ր���3 z�1����d"�~�/�ڊ}�Wc�"CPڨ]��>��q=���Y���nA��yl!ߚ�k���}O�ɢ�c� ��v^Lٳ�7�e��ʾ��k���I��T}����je���P�P=�J��w@᷋�5Fpj��گZ֖Z�����q��Nn�jR��(R3K����8N��"�ntD-,Qb��6�ʷ�8�X�^�:��!-�';�����0�)�n2I���|�@EwN�!�co�ڝ�T,���mTW}B�� |�&Y/�+�z�֤�T���Rlwg�̶��W)Z;Y�nT�͌�;�!8�9��Y=�='��%'�qI^�X�So�k��Պ�FB��K�o���%����f�r݋��D��̼�����	d��
����R%_z
)�{�$9���{K�)�ɹ�8�����e�L �k%�������`����S/�өZ����uH��Knbc�"�7������t���ѐ��Nun���g�˽�Ah���^�by���5���19���`ߚ����Y�DD�Jb&k�U�B���8~�Vh��2d8OZ[�����?<a���x���:s�R�D��'�uN#�k	����?����b]N�­|R��������{��m��d�^C�05MOW�iI4�a)OC�\���:����w�Y�8a���u����}S�?�|X�H�(I4�}���'4��re��]���pV�ԣwԃPp�a�B���CUl�w\�������F&anT�]��4(AU�Ȣط��A�(N��lrZ�٬�.5�FD��S��f��2`끱P�oŝ�m�}+xi3͞_3k�2��.�>Y���Kŕ:�~�W���3	���a�ԧ�
�*k�r���WR���,\'{}�ϗpϴ����/j�^v��?|׫5A>n�KU�B���o,tj/��;���=
oV9�mޓ\����kt-S���P�k���s�Cg\9��Q�j�nl	-�춲BI�����W!�k�-�����Yp[�Q8���xU/�����͞
�l"��ݮL�D��,�X%��#���B�����g<��g�ጝV���M�)Tcn��Xy�^�-*X���dծ��]��^ط��� t`O���k)�5��B�5��M����ɵ�����7���bT��S���� `��J0]�P�P0�����P��/u��OOVu.�{��j��r��,F���\��6!!*��܎N�����$�{\��ب��<�I߿���'���|�kѯ"����q��:.����=�o=�]FF�nR��e`1,�y�s> �.��sb?l�tn5TP�[�^�䉃W��S:�����J�+4�o���{�&Y;���  ��k��s{��M�����_�y=�t��*�Q�>8w�w�QI��\ց(��@��y�R�z�MJ3���?��%)k�^^�U�$�i���l�A�	�r�� e���nC��|qX|&y�C=̅q|��3	�Km�E2�B��5W������I�͡@6�f�B��SX��}�QT�s�#��v±�¡�q���a�	�.�%]J�u�>�ì@m�_ÿ&+&Bͱ���'��[���
�Z�Z9�)����
7�*r�׼TŶP֠�7�*���I#ب%:����pm��ހJ�}N���U�.��u�^;�o��K�,~-��F��~�S��QgqN7\M΅g0g��������K�F�ل��%=[GA�b��_��15�R���/	���ڗ�"P�1�����@ �ș���%L��M�Sy��br<#5U��7E<^�n}ۀ�(�[#g�:�J_u#�p%xj:�"��.�"3��UL�B@׊Ӻ8U���tk>����nb/�5��|zKF�x;9�T���r�H!l,������e��4�/����o3�@0HK�CK���.X?]5`���l&��BB��(���������9٭\��,ӭb�_���%|ZA�I�ĶrR͖7s��Eҁ7`����^F3�ŏ�:�{4?��L"����L��Ǵe�|l;LB!"�"�>,�w� 2F�l��I�3�B�E�7P��n�7-v��!����];����p� ��pesG"�qv��)Q�����h�U
�!F΃M'�Z���)�Y�{!���C�>�����W�qh���Fڀ���=�[*�D����o�Z�`���c>�ȱ(g�܁_]�8��9r:�XU�zw�d�3�ݢ��6��~dDP!qش� D�q�K���#q��������^��-v�8B �6kPt�xT��T����N�
�7][�(�g�U/<h�5Ƭ��;�׬"�G�� �=�M��������I�iO���u�]��>����"���#M�Ix�|6�v��@A$����
y]Ie���^��I�C�j�˭ŏ���"Z{�ް'��һvΓwn��ka<�t���t�=�?��m���7h%�B��D��3R�Z!#v�nS���U:}X����y�{5>K!�U�)�����yYI˳,Q<2:|�	��0����w8Υ�/��.b����Y 3}�A���C�`����t�����S��W~�����;��_��r�87�#(rFxj��ĺqE3և�B�wʘm0������O:��:ǖ����z2O)E��N�� ��r?�;����n�fT��l*{�w�$�*�GSV=֦/d~t�A�E��T�q U���Q��Wϒ������>L��f�b:���(���y��g^����'���T���i����oN96�
OPR��
���b�>E��>z0�g�����S�|(B��տT�?3��s_���>��Y���O��?��900��[Leש���� �����#X�J����Ϊ�4��1�5�q����բ�����}z@v��u����@M����KC�=�����Y��J����`��It��)�sCzNvQ�*2}�scttT�>M��p��j뚤�TU�ߕ�F����o
/���V�N�4'������ȵ����U�P�;���'x�E�OO���IX/�}d�-q.�hBB����|���-t+2�ĭ�i.�=�L�!�# ��Q-�<�ޏ��(q�0(�γ�th��*�ʫ�ST崚�6���M�Hb��'�'��q�g!:�y�8+�g,: +`&�r�Y�d'f2�O�Sf�"ѳyZ��� t��@�'��d����RQlv�S����-���7-�++Q*S(�?��n��v�	��Ýo��*$(֯��?Z�Փ�5KZh�o���k�@	��i���~���6g_��3�8�}����×��f��8�a�,b[�'m]<�M�w����a-�%`z���0,\��;6���n�梻��YS}
{�t���NAי_}Ē�j������B�^�}&�b)�G4}V}W�6(� l1c/��{����X�מHP:��M�A}�����{��@RX&��B�~2�-�Ǥ쐒f�y��Q(DZ���o�z��5K�)^��\_�uߤ�sA��v��#�| R���w%XD� d������D�:s��?=��=��N��/w��O�39�9�+�l`v���p��1e[��h��"��@#��Z�ow/*�G� �^�0KKE���w��ޮ�ٿ���yO��V�Ǌ����/Ҍ�L*:7��{�O�8�Z�nR�������.Vb�o�pm�UU�b�sd*܂�ސk�/i�2��e
}&���I���y�u�zY�VB��������f-�6V��Hq�!��X�����p�N�Ƚ��cP��+�0��&E:��(�~��ƍ�Z�E6x,o��{�H�cI}^�Lx�̿��"��,���la6���"�c��㝃ݞb�i�!(x� �N�69w��a��!�z����8w�k�dj�D�걗Ì�-�h��?R11EeWX(�5n�^;���sfR 0��ؘ".N�Ȉ\���[�u��@���xv��'�[��&�u�IK0b  <���X�蚘�u8�{�,�:s�0v����v^�a�
��h�4�}� �,�Y���"Z�"Z�7��Ӹ��ru<?��uX+��_�m���ԟ{�
׍ c#{�ގ���z����:`��+���*D5EwKqXQ9���\�Q�pWr�Y{Όg���F#�����|����9y�j�X���D3m�1���";�U�J0ݸ���*G���&,���x'y��V�`����_���S�q��e���F��Z����m��:���#�q�C�F���}Z_f���:��B��xw��)c�'��%��+!�<:%��񹡊�lW�4Q��U�k+u�Pמ�z�X.[�j{�vv��"�&-\��]q�`���]w9;�^�?���h�]�W���oc�kV���}���T]-"�dQ��8y�$+�1�/S�g�����S`�je�<d���G������QGu�Ƃ\~9�}r��"����PW�1wVE]��*���� ���x�1����S}�+�l�wC!c�p���s%�`����JY}�*����D4r|�a}4]�X����!��}�)���ȸ�<''��5�u��m-@��!%γ*�B$�Y�a��nH9э��p�Ϗ��gf.�����@넅�Zj��Y��D��t����b��J�̽:�����s�㯛Πq��"�q_����$Y+=w�~�Ϩ@r��{�U=�����PO����K��U�����i,�@��86�c��hMW�y�-O��J��d�L+��%�_ސ�n�x>�mjJqǘ/�7��ݮ؏j*Ї��{�'{;X�5���q�m�K놸I���ߺ�2��5<���_�L�k>m�,�m��j��	|2Ρ����\�s�^J�L��0*{�S�ޝ������0����Iá�s��>g�e�����c+������$�[�H��p�h�P8Uh|��M޿�/_�?@��_"�� ����~�ڵ��u���4>��X��)�7��2���Y
>L�u@�^���|ƹis0��81�a�;xM�g���D��oV�@�Z��O�k�dE��Z����%���?�d������0sDG�^]�t�͐h����fɵ� É�A0J��ri{������'����K2��lې��T�=(e� ��o6�Us��[��j\�� �:!Z��T�2���=%�"�ٯ��/L7A Ђ���|���nq�lѐj�v@��Z���Za(��s�RZ�gޤ�R}�A=�M�^�<cd�-��Y�\�7��{{�
;<���������u} ���Kz]7Hl��-U��z1h������&1w�5�*t^R�R��;8�6���8O]$�ʖ���R,�B����э�o��ص�L٫V����o�o����H�V
;�B�D���V��B�#�r�=;��G�C�ٝ���	���L�{7���b3�2����Y~�?ud�H[�Pk��oU����������npU㪔���O�_������Z�\_�Hy/�m�'�S���w[�~��*NMd���f�'}�;`=��i�O��D���3; ��]�>��@�{.br������Dް�*�:��%~C�U�a�U�'h����&}���X0K�b���	/C�a�Z�ԑ����!�B�K����6Y�n�5�7�h��J{k�D��p0e�?���vYA�%���ӎs����+J�4�"�/4��@�2*:��#�6=���I�WI`�}��g3x!�V���Pb(��?��8����42+߃�`MR�� �kNw�,݄��ZHzoÒ��VGy?�ey�7(�=�.r���W�OIe���J㧐�+��{ m�w�v�n��Q�V
�S��*ٖ������^3(���(](�]�;�������3��N\EU)���gW�����g��=DV{*���d����zI�e�6���,�4��e Tֹ��qn���G�˛��*��*�|ͻ�3y�4*;�tq��Z�.�-�Ѝ�r1�z_3��R#bow�e8;�~b�H{}"���zx�}frn��d�9��sϬ��Z�(Vd�B��(��a��*7���El�5��k���#��M�Z�	�G<�kf{&q"��7O�(�WO_���FZr.2�?�$+����yM$5R|�Φ.�:�TP�[Ũ/�F���
��~v�I���
� � &�+_n���:�2�1Z<�*�h�J��c>Dd�~9�~�Hge):޻Ĉ1(,۬�<u�P�D򼏥|��ִ�K���E9I9_�o]���-���c^�<����L%��l}ڀ�\*�;X��<3D�#t�]^C��6E� ݤ�b�ö^P�PE?�D��GZ�b\�^����9��7P�暨K�9������,���.��β��9���̓�z�]�ݽ�m��Uf�Y��4��̞��z�|d��/a���=pgяiKڱ���Iz4��@fJ;cV}�(C�3��P*Wun+��1�xL�L����2.��y�(?��g�HK�~�Y
Fo��� ����J���>2`���_����߀�S�}�J���B�7��Ѓ%�Ui���:L�A͉���=�ߌaW6�8�E�3���&mV_(���
��}bL�`sw��.ם��89G��k��D� ��ð�����;d�9�lo_����l�b6�s��x}�J欠�������� �j��'�Ѩ�������o_6�PA�0�+Ч�!æ��=D�w���'S�;���䜐z��R��	� ��Xt���7�U�L�ޔZP�XS�x�:�D��Io9�뮼��
�^���3Vzi��Mb��@b�e��2�;�Kׂ<�۾^�6wtn=6~!�E�m���Rx��`�l�v��<�@������c�xh����6 �V��8��c ~E����;��7<�]`�;Ys:�_��+.-Rr�������S���#r��R�W��4�����3	MH��=[;}��4#i�,Y _:��7��;�;�Z�U_�^'1�G%��?�Cк�>|�e�Ξ=�n�=��	ZuR!�7�>��h��ϊ� �_��QSW"2��߫E�Ջ������h��X�	ԙ�*@}�
��ߣ���I�&�=W"��s�����VD�B���xҪ]d�5�n�n�<-90�T���$�E�g�@�L6zUۡ���.nrw�jd?���'�~�<����r��Z�n��)i����q��}7�=vˉ�� ����2��(�QK&��t���G��̈́n_G���i ��"�f-!s�o"z�(�f��*�ؗ�L����e����w�h�<{nwݬa��R�B����B�P��zIc�:.�"�U�N�{�j1�:��s��g���)(۩�ȋ}^�+��0�h�e�!�Ȉ]���;�qeJ0t��k g���>"F�1�n8�s>@X-�3�*��?F�^�S���g|y�@�JjT����WZ�4�d ����'�tgy�B�P�F�3�&�����O�|�]|b�
{�^��] ���
��^I?>a�!S+(��ߗ�W�����Ql�:U�1����A{l��/ǿ{,�/ȅ��8s2�6���8<O��&��������Un�W��:%�G���NB	�L�E�j�4`�Yd�C}Rrs�J;��mBB���*еa����_� uE�9Bʭ�m;�Ĩ�*v��%�{���y����q�Y��D~f����}���!O"�O2#@�Ű�7]���P��Lg�:�Ӟ.����-翹O�5�����P��C�����]S5��.O������i<R��'�v���RuD~�2@�h&��+����[6۸����.�	+�BL��{����P�K�4��3�0�o~2Jn�޲nӿ^�^5�;E�㍛��!��z�}��<�z�����E>z�X�3�Rw�[V����P� ł�����/6?�P\�;�}..�HH�,�/&5m;�$X�W�={yib�i��}|�{%veH��]�ݲ2nu�V}ƶC��;�S5j�,2 PƮ
kѸ`ٕ�d@�?{�C��U��n���*��K'�8]/�#�����68�#�����{[9`���뛇D*BF�m*�0#A}��Ȕ�6�|݇��gV�@�����h�U�@Q��U��E��SF�
�}�[�\�����b���H��+k��C�ތ��,�٧A�&M)U�BO%�N���`��y�g���Hϖr�C���/��Z?氪9F�<ԜOr�(�W3�� �M�ǚ\���6��)��N�w_�gv���N4��5��W��_�CE|Z�}�'�U��G���2U�K����qn�����P����!�.�ڊ ��ݮ�J8;��A��5S궻���#,� 㥉���m�9Vk��N�ǹa���}Pdԩ��ln�����aӯ����N��̾8��� ��t�	H��È\�\k>�&���yB�:��ɨ#�}k�z�ǭ\<��w�F}7D�)�0J��Cp��#5'�m�&Q�Sne ��|pP����0Q�#�Wq��Y�֘����v�.@���uYf	��7y�!2^�F��\�XP���i�FhG��݊�YU�����ȭQ�o�)���0��it���o���^7��>�,Y�I�]�����l��+ƺ�^Z��T��;�(�[E�E�E��tEbW�O�;��s��"}���ĸ�Op��~�f�q�X=7It]�:=-`�� �F*�]#�nVǋ��$	`jq9�Ւ�n�c����"9�x���:"��a]�V��HGQЍA��KM5S���Ң�J?�>�;�ۓE˩Hf��v���-3��=rH�f�A��������&U/�o%t�[�&b�O�w�Ȟ����m}��)�sx@��+���:��%���R�AN����"����V`��x�ũ��5QƄwt�L�w�#7����;�5D	���a��S�oՔ��غ$W9b�?�����	�C1X�+M8��8���7k�� �H%��۱��ط�Ϸ�Ռ4
5�3դU`��H�y���wz@�wy�-_�"9,�qg�6�,�c��Y�e�7����r�ߝ~�޾U{d��V��7� 2v�J��ps�� ���_S ex}��4�����Ϫ� �'��ZT�c�#�ݎ�P��6���?��$�؀[��5���E�Lz��3� mv�X���N���r������Փz1V}x�ϗ5�����O�X���I���lJ���g�K���D��m�/�t���²�fr�ŮF�/|}��ȳ�	MB�vU���'�߄���7DZ/��}�B|�2���ŭY�.o>�������'`Z��e�oF�?�VX�k���y�?�4y:K�����q@��ߨ.�}1�v�d��Sn���g����y&I�����e'>���Q�X�R\f�\��pc9w���70��ނ��\G��������y1�Z*�Xv���f#��gv����M�,�Vz�f���8���&�9�4rr������9�vP����Ι������դ�Ql?Y>|��������0L釤I8N=nO;v�<��ư �"SR�8)EY�P1|`Y�ڬ���N����'�aQ���
lI�V��d�E|z"�P��DR����\{]���{C�����	j���;�yt�5�h�v]S���N����{��6����T�fA�v����"�����&|k�9�#[�`8���A?E�$M���<^}]HV�r�i�d�:�����F�K��q��_�_3�9~-��̩��}8�ԺL#�kW��=���[k�_����S���=k�Fc�d6���L��D8 �-��TI%b+�o�?If��#�R���ud��U,6�P���P}fƃ���-@4�GV�S��=�OjHTa��.��&�K��~äp�خ��-����tF�6$V�g!��ݨ�.��H��i���{����m.��j3<��h�/1'쯍�"v���x���7��4�D��^����-2���5�N5�h("-���(�y��%��z3֒r�豩�.�Y}�M� �j>})���qU/\�'<��cx�5�!�4���i�R;V�dTz6��!s�]�������ϼ�p��MפlA��H�����([Y�5M��h��&��9�W�ߦ8�v��%�U��+57�A�p�����pi��t�����ĺ_�t��=�R��@���tAE�r096.]�@+�>ԕ���}���q?iJ^���a�i�[>��LR#����OE9K�쪶��gfå_D0F���,A���[v����2�vZE�C� �9��E���1nC�d�M�+��p5���}I��c	UJy�H�[q���?DMѻ&�^%z�kH�N�=/|�A�W�S:�W���ؗ^T���-)�쪑j	����|w���������/hr*^�dev$&��~U���\$���'�w7�jT���_y����0a�+���3#�Ԁ�?$N�7h'�˲��T� Ҥ~�k�fVl�+!�hm���F����{*�*�����K�S�ڌ����K ���W\�>M��z��!��Q�葝)YO�\�Ϲ��@�@��w����Ǫ��O��J�%��$�5��ׄ�����-�4����[�з��R4Y�&�MDҙS�X���^Fݔ!DN���/�_M_�:�8>?0��K��*bvKLHD�t�F���-���E�?2�{�i�������������S�:��-~�em��Pd�޴�e����nbI~�ͣ��I<�|&��O����_��(�_o�933�����=�bL�ݹ�O�$��s��mnv��2 ���`��O��^�0Lm��_�y���q�Y=e>}ܝ���O���^�&�m�+!�h�Ͽ��o�Gby3�U4Q8�FHU�aq�|ʧ��?=ޜ�?�Ej����ܒur��c~��W-�l��w��PQ��'n[SJ��!���5.�S~j��o=���{�ɷH���y<������ǣd�m,Ϸ�]�����M�����߽0-�(�v�v�%�=mʹ�ȏ��Z[�<h�z?檕M�ѣ��ߴS.̷��1ſ	 k�<���-�����K��~�w���_��{���fkv�B�>V�cd	$�U��}A?�~���>~��B7��|۲���~O��Q?ʢ��hB�V1��2;L�F"��?>�ݛl�����J��\��5���Գ��,��id%=)�X���j��}�s���	� �J�3�W
���%K���e��Ok�O��{'�:�*6��,�f�jP��js�Qo��Z���b��[��(<�t}���s��o����Ío�tzM5��KL����~�����|/��{��7���`o�$1<oc��V<k��K���]���a�JV��G�m�&���@
~q����%F8��ޓ�O�g޲�p�穈]����	�u�=�QĀ#��}�Ҽ�B�#3����u�SX��ep>�d�8�g���]G��.ć?��sj��a}�c��G=i��5jK�a�]9���%:�R5�����r��ؿ��R2�q����Z���ꁓ��9�5�j�}�i��'���+{TA�o�9��!��������᧙$�j����o�f�D֢�nE#����o��/��Ņ�B���3/ǘ����:��C�V���C_W{��K���t���9�u佨\�;J�;��k8823�(ϙ~,��6�n(���U�q,=�3:�C�0�4�I��г7�ƂP^�K���\/\�	p���'�.����PQ�����HQ�ʰhQ�<�q'��xCܵ��݉-u���M���}2�ݼ?L	�M��Q�-3�7sL��G��n��1�JνN�.�{m�!o.�d�3EE5=����r�)x��^�=���;9�7���cuܾͧ7r�_W+X�=Si������|޻!��<nOT�����#%��I9!�ܶ��\���2x�q�K]����r������{t{��.��-����,��ɹ������|��?'�C�[����c�T��D�!w^u�PH��V������Q�\��sי-;�C��� ��),��EG�n�W��گK�ː�;)n}��o^_K7����{5p���7�u��QnN���.�wlv���l�fR�Q�z.��6���/���� �����0;'w%97ћ�q.DĚ��L춾 *�Zvһ�`c����勡|i[�tC�ڄ��陙�E���f��5��Q>֣�'Jj���NT�^����=�iJ��6���V|�Ac��6���g�qҵ���N�Ǔ���$���4%fmY浌��m	��G�gI.�NCE���<7G�$�v�?�\�^��==2B/y���G�>��i�a.#�7ս�
e�yt���?�1���p��k�)��o��g�)���1����{�Nc;NP%�h锷?�d.nb4S�e�����L���-\��M�`s�G���Ӌ����š���ny��ٛ�_qLi�ſ��b�Z>�� ̂�l�|�E�>Ϣ��D���BO��S^>6����I׃���o�<�U.�F�,`B�j����o�u9�����y-���噇<���4��a!����n������k��.��BFeS}�K�~����SC,.Jk���?�s�z�'�ְक़��e�
��SG+�K/FW�d��V�*Ķ��Z�{��䔽�uG��s7��W��D���L*G'7Az�Jn��Z�б���^֮y��=���`^�b�y���i_���E6~�̔=�����m�	�J΍�i݄��9��Y� ��ǎ̯�bN#�P}�:���ot�2m|׻VC���(����=��vn��t��&ԗ���V�7-`����7�������W@E�>�()� Hw�* �H��tw�����t��H��"ݹ�ҹKw�.����{\Ϟ=.wfޙ�yf��{3藄����l�I>���k[i��f;#�H����� �M�
G��!��h�?��j�*](�ۻ����_.�Z��沊4�:��&@����I�f)(�r �����҂U֌�\�]��;��k� �$�l��|�O˖(�^|z��Il$K����1_?�.eXȆI��+RH�Ҙж~�7)�t�6F�`�:�����Q͇���en[ba?�ʡ��>�GW_�����d��/�H�[׋	zN�Ҥ�OC��P�&��'M��\6���B�Bkc�;Kq�,����<�Ϻ���`�w�%�ц�h��Nٟ-1�7��ۍ�cͻ�v~ 9�P��8�i'ñ����̟U��\�"�OJ�r�br�m��ߖG�E�6� ��J��7�.�s��*�"VJ��5����hRf��z�k�������T#�C��s��&�^���?(#/c���1���+��6��!ls���-���]��i��������ܚ��#�;uV��k2��Դ����u(�
�[˵����ǶX��muD���S��rT�5�w�ѩ��L�0�;�y�ʟ\�6d�X���-��"wm�G�1/�g�gZp�d�*a1����t�k�m�K����ɹ����5ҿx%�F�z������y�l�a�8�A�M˿	�#�9Ҋ׿g�E+��ϊ���(슰�.�7�_�.9��������䮳i��?j�Q)��+�����6iu&OP`�F6A��Ɣ[F���O=jϛ�3�;�oz6�?��Ǉ����ga�
�nP���0�y#�sC���ʅ��Ͽ3��|�%�O^��H�K�$���"�d��?��Ѷ1(ߤ	E��|>�����q�卟-}랖���?���D�V1e�˻��d���٘�-eQ��7�)�QT�p�|��節��,�$�:��
�e��盧Y;{y#ǐ]�Q��̼a�]�`cVxZ���X�������Q�f���B������c��Nm��؅����`Q���i.T�iԄ��RD���}���Aر� ����I�tr7��R#y��g4\~�i���D��`H�l�2�Js�T�#c5�W�Oٴ�� .X*��Ao^�M��P���Q�f~ �N��z�� S�v���6��0.��~u*o�Y�?�H���ʪF���=tJ_����_L���v�'4	�-���^]�É�
z�RH�=�;�����e�#�?�l��C�U����n��6�e��	7�'�԰�3���{"m�u���c�j^>Ѵ�=������j�kY�7
�qn{C
�7F�歶ܶ���{l��CyU�@?A跆�
*ie�-���#07�^e���N���<JT!ɘ��`Jȫ"���	��aB2)�!��Q_�qS�_��a����F���ב!bA���qWʷF,��=w��jv����[*�a��g�':���ה�����W,`#�ِz�����A���J��u��dw� ���ꚟ��|?RQ��iop%�X��P'��L�k7STA�S�͵��m�uaWY��ʥ�")u2�ה# �O"3漈��Ǖm( �=��w'�(�A���쐌��D:�?���D�Ġ�� �eEo��Q�x�.�4e�0�DK$$�c�d�5c��f8���(MS��l9��l>H��s9WjB^��A���DA��*i!�v�o��[#V�et��_�:���{հ�~u�#�xy��j+�����󧊐�����q����r.�1kP\8���m�T]\,HM\�ȷ�brE�+&W��3?&��G��Q��7&���˗O't]k��1����,o�*5��P�?��c*��/���WZJ/rlTu����%�r��E�o����Hh����1��?[��j����)��+�� �K��aO<�j�����;���Oi7M�A���h���|��a.�MTh��PjL�q�D|n���%�u�Z�>�����6�v��>2������ířJYt^�x,�(��kF� �S�@6�F��X{	Ɯ�4��3�	��{���8� X�S����2�!X�򊆳����G`*��ZqzO*�v�"��:\}�g ց����ö�p��Q��0�+eU�(B_�N�&4�XU�y���	E�!~0m�v��U��Eq���"�oó�=��W%�a�w���*T�;(Q�1�d邭wG�B/�7������.w9�G��|e�Wk2�*�UƷs�h��y�BA׭7�C{��aI�yQ��e��[ŗ�3�7?�ݟ��npS�8K�nVD����GT�薉W�C���[?��I/9w����Xj��76�PVR�YA*�;H������Mp���9iЮv��z�Q��5/ؙ�Z���L� ���Pk��#� �� [%��d6K�?�]��v�l��7���t� ��߷g���
ǁEѸ´�}1�����(��)5a|�;���8N[q��u�0��S�0R|/{��i�ԃBWH��OҦ:�q��Z1t�i{(�
�զs��~�5=��1�lG�!��-eu�+sb�A@#�k��iL�V��P�Wa������J�k�}�e���6Y'��T\�	&4�������ņ:��agջ�|��� ���v�l���?UU�Hؔ|!�])���l:���M�yIϩ�F�������
!K��{�" �
)E�"�+�I3 �+&f�S.�
�m+��n����CQzC�dc��ݟ�w�f�m���8��,�v�	cӐ^/�NZ�sL(�����~��!�N[��H�llC��ݟ��A*���S�^����3��ʜ���
1k�����~˛H�ˮ��J l�e��l?���x wX)���\��}n�+��x܄/-M��k�o�����U���AB�V���LG5�9άՕ\ <�*����XX+%a�Y��ks��ek�\��G6 :M��!�d��1֗����i{CV9�'p롕}��"�w_�-9K&�]!vj��o3�`��|�yA��ђ�_ '��kL��l�ai�k�����M���x�� ��؜jVc�������I�մ�!�Y��̏X�W_��#��T���W�8#�g��~�-T���;�L��-�[�P{��#]�`#�N��(��S75���a�3��j{�ʝ�V(�lE#Iw�M��RQ��b���5�r��9��ǃ���grM?AR5���R�4߾��=P:Z��f/������~�zM�N�4��N�Z��'��a�>VY�K�7���vUCM���Y�t0A����}�3XPy
���Jy�l;�xAo��w��U�ɓC^�/�q/��3��X��r��ߞ5C�gy
���)��h3�å3UP��׭��!��6G)"6�]�2'�:��j�Fk@��ބ�0�p����#�ڒ�19��V6������Kp��U@v�4o���tP��Y����nlZ�>"��`y�3`[��������Y�0���ͺ�U��6��*=ɉV%�X�3���ݏ�S�ӶLJ�69�Bx��;�����_P�F-�VT��#\�z��W�b��@*x~�`��v'?\�oVc���2��Ό`m���j��t@��>=�Y�p�E�f5W��*3+E`�`8������*�����D�[pt�~P��d����!�Q#�98xQ`�K�>ʼ�����ߒ��݃^Rj�]��^o�����S<=�Czogy&�&��Lp���4nX,3���࠾"T�HѰ��"6���C��o��2�~�Ӄ\;�!r��ԿȌY~�z�BEW��]]E�׾/�]J8�)ֲ�X��sǉk���;�"�.�$�层��1Ȋ��|��d�Sʾ��2�&�V��{E�#_�^�{�B_�S�4����R��i�v�+�4�u�|>%ew��vI�d�~�e
�`���q�!;�g�횼۠����I�/L�+�����|[�*Nnl��O��G��FFVg����fZ��a�������amk�,����0��aJ�bN�� ︾��m��d�I]=��9����}�і<���Q�V������:"��n[SQ���O�7<�E�	kYgbp� Y�v�h���o�@<�+����>���Q5��]_��x�������fW�n�N��~�Wv��¹^6&Yz����~�U�@a��v�igr���~=c�\ o�S�-2갛0i}�6�}���^9��ix?mÒ��F��;ҷ�V/��P�;GA����)
k�ڮ /���?Lc�����ŧWs��z{�����(a�1�t!�Xҧ�����[�H����&�|���F���	�e�<uȳ.�U?��a
|٫�"ET��5l�v�e{���yuѵJ��¾S�vUv��d�%`])9?���`�_��Ī�<�_��Q6a(��Z����kv��Z���Ú� 8Y=w��6+��I�Q[K����.pQ�9j2>wþ4.}�J=��w#K�r3V{� �j�wJ%����JH�AA	�M��P��K��c�+�ZK��c��?+���.[,�n�2.�䩿����a��^���O���4�f�5=ŵ,s��
�~��ߤ�/�'BO	*N�����j�E:�S����P�����31�Y�������C����B�n�Ϊ�������jMӇSA�o��c�$	_���*�:�O_�7"moRl//���=][BW������D���(|��1YՂ��~i�/���|�%��8��91-L��=ۻ�Т���c7��gƬ������1�S�e�r�/P��רo���Uf�����(t�ޭh�C׳�$#�Ѱ�s�Ym���vR����1���Į�#�{����4���&O��V$~� ��Q�躤���[������*U�Mh��b���Ě;�Ov��!?��E��D�$��q�n�7����K���6�@�$Ӂ[A����^����Rjo�7�3;�a$i\�?J���o#ѻY`���';B!��C���� �D� &r�i�mky�M��/qOL�P�B��Q�8j�����X�7��/$rA��;�sƙ��}4_�^HL�"������n�)O>5�9'�?2�=lE�^����e�.��#(�5�����
������d�=ˀ�xnu�	T!foRS\�2�E ���U��op2����%4��O�B�lu���u�QY��]�yyh4� ��y��Vn��!$)�+R��Hа!��J3�������/7�n��P���#���I��U����'3np�e���ee��_3�$�0�YYU9��JCwR�y��⼑�q�l��Aj�h�ġ��k�R�q=͐��( -X�z��$���\/�MT�|�>�����郦s����1h���'�P&����f���ͩ��G�MDH&����'5ݱI���ׂ?_�B��C>�&���܍�%�1v�(l~x��7ғ����ک���{�u���W�l��KH�8��ʈ�e#�ÚL$ݿ-���~z8vp㷝vEY������.��ɕ|2���w< �4��ð���XH���pZZ�8m-I�ņ��_�KK���OU�8��[/�IEɋ�(
4�z~p�3��˼��B<! /�9rN��83^SE����'p��C{��4�����Fn Ȍ6�~�w���s���%Ue����(���U�?+n�~�y7�D�U*B�` �΍f�-R�"(������+����[{m�q&'�w��ZE���'3|U��6H�����9�|RT#��dP�ɖT��6ݧ� y�lGt*S*���4��2�DH}�sחH�
����������Q�j ����d��ggeu2��C�7��Su��>�7��EF*��%/9�.�V�q�NJX1l>>�U�� |E�V���g�Ƌ�/�;�қ0#���ݜƝT�νG۩C"L���8�dv:���R��
����߭X����M�"�Z�Y�>VV	i�]��g�G8�Y��gGF-zu��(�2��x�I����q��.m<����	�b����V��|f��&,��07:������G���0 ̯��OI!�C�6�2��}o������OI~��(�./v&��t���p��9�ý�ܬ�H9;I�Vp��Ċ@UN����(R�L����� Zr=���Rr��^���ǌr�1�h������7�5�;3��3+�d��R��,�7��W��燫��s9 )nW�Vr����^W��`u�
��B�֔/��0��7b3��*�,@t�|���nv}/���ۙ�% �Ʈ
ɓ�&7ަ�㈌E��3�FEW��d������X��*ŏ��}< v]B��L�����m�i>�l[���.�(�#���`$�~�����>��gf��$U�� ^� ��0�z\���)�1�P�<%�'-a����o&Vi�-дI���S5Q��ɛ[�}���GSM41��֟�-h�%X�MD��.IkW�Z�U�ɦ��2>�4.��8M������I1�D �[�H/�fCMJ��O"�<F��+7F��b�0ܺ�G0'��$�$�9*ȉ�U�rہ�d�xe��)�JI{ח�h�,6����L;��d�2= �������;Ԝ�&z�V����m�$���e�Cu8{�Rϻ<�+7'��Lš�8�����nc���������g��b��^Qd�4���V��B����$�@���k��ldȢ���7Կ:�ԦS�pv����r��jh�_O���������aWr��!Es"T��/[S�?Y��(��QF����h�{������:Hm��y%"�_+f믻�}����L>%�3�)�=�Bϲ�=�1v%1���ۑ�i�/wo�#��;�U_yh�|�y�_h�����S� ���J���bp��(ҹ̣�U*������Y�ն��1|������g�G1����/fuHv<�H����(3HI|���ژ�m�����t�cZ��2(c�[��7��cy���R��o	�&��Ƽ!��B���.f��~��
+(ޠ�%N6�@K�z6�y���6m+��"�C�A8�{���%��𳎛b-R�K ��ѻ��*���j�H5�\�4�K`y�X��3<g��!7UD�_n��w���~�vwY��G�	��?�q�ʏ~<�6dŋ��:K+�1����F�Z��ܯ��
��2,z&;'�r�\�EX�4�U�Φ=t�~ػs�n�R�����jI��/�
ԪE��]�~�)��‖�G?LW^z[~��Vu�z�
#v3��d���Z�U[���M��MWa<e3L�p�c��du��&��
����߳����*R�[�4�&�ƨ�����ch���ά�<����M�M. l&��7^�ͤ�ռ�f��CYQ�m�ҷ���%��?�4��~�w�@a�"ax0A� ��XL#����1��:�Tb��WC��g���@�y����I��d]Q!7��S�����jW&cV��?�NJ�ny})���ēP�D���5��M��Wg������ٳO��C�n���m7�B@X|'���}3�QZ�@H��],>�3֖�͝���*�&���������h���d� ��ï���"�G����Ы��v�fw7z���`DZ�WÈ��%:��Ȳ_��c����DQ.����rD���"/���'�0sl2����������ag�ДW��,&�d4���g��Pc�w�K��=�xy:�8̓uZ�&���[*�
����-�H�����՞wGa��'�"ހt�������=��#N�nY��æv�ew�羛Ԉ3An�&;j��G����IC�,��4��"�ע��^�k�@��Kܗ�k��Sl��B��e6�H"~O��2㇖b@l^���c�9+F.��~�MoI��AH��~J��t~<�q���ny�s���m[�X Dl�������]�OCb�Cv��{��{���M&����U�k�2=����k�_�N�cv�ǣr�y�g�Vp�҇,��ry�B��0\�>�[9�~�P���4F7��ɿ�|���M]Z��r�[� ��;�7Ïi�6��ae�=�3�)�ݦ�Ϫ%VK0��XEhK�o���+�2a��=���{ըĲ�z(Rf�Aƒ"HXm�^�w,�L�jA�qg�q}W��O"_��5�~,�@�-I7�i�ԁ��B�I%M�g�\A�k�x��aD�Eȳ��|�~��8I��e}�n�t�hb?k�[��u
���\�-��A$=�eۗf5��=;�Ƌ8�y"Gmj�#$�S�tP{�����]l�<�������Y��':��A��1�O�~^�6c�uu������$`tl �axx��m�Y8�ħ�R�I�vg�Y�k;����P1k��:˴%�"ѳ�?K�������6�~@�R�*0���M������j-ֳ�BV���^|>�V���5|T,�OQ�Q;�t��Z���0��ę]�y;7>e��E�]��C�4tG�
'��I7����Si��Z{��l��\:�o�+�C�v��]��5)����nG&Mo^��;��&'"��_ \��Q�O�Vv"��l��8zx�=�����;cLn�ko�~�!a��A���8��7�@}�g4�\�3�,b�J;��4F��<�<S��{]-!a�>pi=|��|Դ�9F�l�5d=U���!T��������~�N,�m�땦���#  ��
�EB�v(���k���P	Y���Z���ɥ�ȉ��3O�d����������+z�D����s���f=��׮_�}��T�zx3Q1��PV����5S� ���Qh��忭P��O���Y�	�b�eR���v�m��9�w�o/��Zz4孩�'��/��hdB�Q^����D'k�h�m\^`�N�4$ o�����u�\�*L�	����Lq����*��8�M�O�E��ۺ�Q����"��qP�W��Y���3��� �A�Kh��m���G�u�ϵR�GĚ�KU��a��!��W�>��'��K���=�i!%�� ����ъ5g-�`�g���sh��1��D~\�r�-ֽfu^����9�W�L(l5ȯDz�é�I/c�E�JFG̕�> ��hK�vK���m�oۢ��\�59h�^Α�1y���IM̿1���96֫ifv{L���Z�
��\��df��g����v�O&�k��'M���ݶХ@)����S	�8�����Lz�G`͢� ?&���� �* �;NB���b��6�J�+�p��n'+�]�q��)��Y�zL������ U����q�a�5$ !�� Q��GX�u�Nq��|O^�Nn)��T�^�����sX�M��{r�rLW�Ӎ�{F�Q�5j�<�����Ƨ���*��]}�<����j�I]�Ѣ��"Wۺ� @�d=~\��8������yz7��'pjt�FV�\�7<�e���-Qw�F�}��_T=̺ۀ�ҙ�ؓ�]{���?��<O,���Ħ�q��0�k���u�:�d��$ۭ=M1� l.�����d�.\���¡��r-��1�~R����$PȻ�z��(JK���ITx���=���(V�OeX��i�_3�⎛�Y�N��MTZ�-P3xr�R�Gvi*|��M	L[lMva�
&{9х�����rv�mp�U��=k�뻐�=E#����e�,K���ϩ���0n���mQ0�����j�М�:�6�����Κ�!a΍ǚ����P���?2���+x��O��+�d��h|X��f~��J���[��9^����Ӵ,��MdL�� B�0pP�PhԀ�S�d?�廡V�`k�i]��`����0��8�<̎钨>x.�@�@�	�нR[�Y���^/�G"�����;N*K�E��Q�&��( �BwR�h�Ģq�5�M3+ �T/�/�1�|� ��wY7�/���'�|�)O��0d�57�$�|��6��� �Nv1/Q��z{6(�bU�a�t�t��Թ���?7+��V�S:�| z�L���������c��4�5�<bۦS�'�d�͘.X�C�dzQ���]�~��+�,�4#U�WnB���&2�<^�'�\�I��_TJ�Dڈ��el�dϦ������$����$PL0�l��	~�T��/���q)p�ϝTl���積�ڳk���	�p�K��ߑ���{���N�N��)+ǟ<M{�<�jDÓ)��k��aO,��X��nE�O6'�t�X���ң#�/���R�F��8]�)�J��['���X)<
��kv�*�z�II7��w�QhNL�h���>@�J�r���y���ſT���+�n�>G��
���=5��h�c�9���1Pr�m�~.�R�-J#I��!+|{�ߌ�6�:�i�ن�p��5��קW\a>�E�'���Q��eŜ�ڋ����K�Q6�\UJ����v����-d}8I���4����c鬕��S�n�Lc�T#�f+nqt�t0Wn�q߼�i$}Cr�'����m8Rh��c
�
�@"!7Xu*h	�D��{yi�J�N���{�v���&�3��K�V����<0�Y�Lr�F�a�Cq�f$M�ӏ���,��ZV�TU*Ƣ[\.�՚�c��ȧT�*f���\��z��1k��d��
�Jj*_��ԛ�
d�d?<�zTP��̎��ke��K]��U�PhN$Tf�m��(|�Z]���XuYQ5�^/�I�jێ��;�l����G���E풌8��XBJ�����"kEj`q�Lp�ߩ�p���bA~bOk}�%���T�3,�o�Ig���g���g�E�����59\����(�9��x_!��^��[h�j��R)<���e�� ߔ~���p뗏�����߮�4��a�:gDh��t��c�����o!�̷���Yܭ�F.��ʙ�W����o�%6q�?���B���u}-�-���a�vz���2K�
5���S�7l�f}df�ݭ�@#ә[�+l4��X��:�1�:<���0��c�7�8��:�]{���I��/^"���Wn����N�r�'JRïg2��Č�L�N[:����$�,7��-�up��Oo���ش�WN��l
7--�^��26|q��L�V�Jq�X<��5S�x�,����Ƞo��3*f�Ә'����ɭjNX�u#!��Sߣi.X���L��+X�ׅ5��t}�к�nV߫�@թ^3���a���B4���'���D��e���ԇ�b�Z��e7�卹5�� ��25&ǂd�P�u��c�?��>�)ɕ�J��`����Q\>�g�{��4��M���o�/&���,o���	i�����K��a�
��_�4[����ܡ�Y��D��,u�m���v�b�K��+`�tb�8���=f=���H5L����0.�0�Ӥ>��	x��/{�Z��L-��n;?���}�p5R��K4��5��b�D��|Zr�t���d�? {!,y<ĉ]OǣKF׭3�xU�HMg)�u��5�ߌ�ף<�e�W�l��cr���
W��@�V7��1y8�,���y��-�����lb��{H��ߌ��Ū=�ȫ1�Zk�$@[��rȊӦ¢��7�t�P��Z�
��r�@΍A�(|���;��C0�&��z��쨻�U�.��$��W�[?�E���z�� ��?�i�K�3�P�'n�_��� ��y���H��6�>�G�)��l�N��0��lX�Pu�d�-Ȓ����A^|��ۺ-E�� ~���Z����L�0�'�X���і1�H�̤�X˶�w��Fک� ��Y�ib4a�7���-���
��g8Z}~)ѝf��e36ב��'���5� ��D���Q�㌍d�V8`����T�Z[�����O2���輪���FM�M�����"�������_g��w��dN�u��P���5{��;׬�Nlvc��@	?���I���.IҶ��%�ra�S��_�v�R�u?�k����ZD��р6��4�y��/W��B2*<��#UsH�5�����fЧ�Y��LIWp��"H'xv�>_�$�n���,l�&������m��v���j3Z80���f�r�ޤ��B_
,6J
������C�����#d�j������ᓕv�	9M �exY0��͜]ޛ����fm�j�IJ�%c@�ӆ>�j�i�7+�^���sx�^�-�G��(�Nk�k��J����x�maT[2)�/w��[��C/vD���^���T�:|4��x��`7�J ����Ym�jAV����C�Ut�T˭e�47���/���[j�-���]W�I,2T��K��L��B�=w9U�d��������L���Bq-�Zב����;��aSq�/>���J?�p��I��4����B#�Iy�'�;{D&@.�'���I:�����c�r�����mְj���6�ǲ�![n�(T�$�
͢OMS�	+R&��䱶�~���^��[����}-���fV���f/�0�뾥�IQdV��|r!ޜ�x~��gO��q9��+Bg­�\Iu�,'�Gw@
ɸ��J�8m���Y����G��'���}he�C��L�C]�.�+�6�
5��`aOv��N���w�7��i6�5���"�sen2�@8&��+�c�L���WueҸ�����7�e��֎�w`L�ơ�\Ԁ�t1W��}�l�"�v�m�:K�y^��2�y��6I_�J�~`��e�lqO9����|]kƁ���Y��.3f�X�m\J��"�0��,`�#�t�ӝ��^�	��5�B�����j�$T�w�����~F�&|	y_�6nm���.� gRszI�� 
��kf�j�>J����­
Qe�Wxh���o��Э��H�Yn�Ꚛ��|_�:?����t�}���|R�d1%�~{1&yZn�G� ��fm�@�͟��<3�U �{��(���h�,�J��1���f��b���\���.��'�����	���cx쌉��a�B���`>��F��`��@��SV1���rq�h
:����Juj���ܯ�т⎔_��y��@o'�@j�p���S�}�w�� �s�Nj؈sn�cƔ�
�v�g��|5F>b����h�,ZY�5Vl��k��|���|���,-�ļi�w;�q�Qf�#���k>�맏��g�2�R�"�g�) ��ّN�w7�����|���#I�$8^�t7���� x������w�N�t��y^�Ӷx����X����۠f�FH�j+��Mr����ß���C�kQ�T`=�?wO���
���}L9Oe�泸0_0��lu��%�������PI�1�n]��s-[ �i��9\jj��^�1�wr{����dPk�!+D���y�zr���+�O|!��&Lq�s�i>�w$Ԛ\z�GY�J�b��G�V6�P�$"{8�Z�P�j5�8:��f�j-K��\�J5�Y�oh 6�m<�s�-�4�r�gϫlg�mО�ScF���M��P��:_�I���L|�)g��7�hw�fsm�u�����s��) �d���S�a�ޥ\����;��J�����I��x����zS�%Ł��I#��)���y>��N���
�N-і}��?�q`"������L�m��f}��1�� Cr�H��}1����������oI�	�W��W�_��~���K��o�j��P֪�pW������F��\�f�_�B]�ܬ�w�Z�T��w��V�=I�^-I,��T��x#�{�q���,�ۻ���K!���_r�׈��$�'7�@�:������0L�	��j_��������"7�sd�Y�h�9�)�� *L�(�(�ON�GO�o��2D��C��;�}ҋ˭�������`֟7!z֕;�T��$Ǚk��f ��!�� W;�߇�u^{j׻�;�d`:^��$�����;<��q���%��c����3�{
�᪣w�bS3&��y�B��;o��^\��եܠ`�6YB��n�_ݖ�ר�8�C<���<�.���)*���咏E�R�A\��T5�L��S	K︕�]:����n���Yg��_�7�٨�!kH���E���L��v�Gd��)i, ��5��1p�֙�Z�%1We�xJP(�NjJ��{nN�Z��ǥ>8��:bg���`&�I!N��Vؤ���pD�[xf|��p��Օo��i�~�����G[L��U|�3���^�`�f�-Ӓ@���N��<�/-t����X�Fs}�/�::�b�n�}�Խ�>�85��tG�c�4�����|٤[j�s� ��۬U᡾,���������1MoNg��'R��/��j�A��ϙ����e���� �ٓ� �O��ɓ�FԷ6{�A�"G���|�g��;Տ�:]؅��/�2$L]#j���<��_OV��.��{����4Go�"�l�$]°Ļh�t@t�����"x	b�w>-���?�i��j,�c"�L�-���`�}\G������a\m��D={��>v���w�H�cTi\�61���{}�.�VR���2M���u/W��l�wl�芛��>:��6zBީQ��l`&-o�e��:����>Cf�*^���2)�\[b�ˉrg�y�0�&��_n�8�5#{���ݶ6>]D"��&۬?�Ť"���ϩ��n'_���{J�#����D<�D$CKnv�s^7(�Ĭ�z���D�t�eD�4n8sc�u�h\����T��(����4��p��cc����S�o	�87�>��ѿ3�*8��4H�=�
�#��p��(��A��.S��y�$d[P1m~�?;�h��B=/�$�Գ)��PH����dr���M&�ՒT�`IB���?�Ȓ;��g���裞6�(o�M����yK�T����Ek|Z��E��w�II�JL�����%T!�I�}ضLS��6gGs���<s��t�L�x杏��n<�?`[s�5Fo��y������-e!Gy)qk����p�L���iJp�"��h��F���ߪ�Z���k��&�T1�٣���t���0�~赜��ǩ����г�
��{�i9
�-��ܳq}�H5���^Ѿ�E��?����o�k��T/�m��Y�^�M~�����Ǘt4�V���;p������ ��ٿ)�*�aZ�w��`1��f+�,�s��0����X���c���C"i=�6��y��b��f��r��J��{S��o��6j�ㆹ@lR$s��tҿE���M�X�$�gr��o�j���n<ˬ�!�F�}t�K��uJD�5������JO���݊��8�kSϚ���/�u�ql[�84�N�f\�]����z=�y�i6:�/�N	r�)P�*��W�	Վ)��u�ΕrJM�Z��3D9�d��5 Xn��ț�$?���u�(���G���AOك��(�lQ�_�]����z�ޜ!P�oS�g�K�����E��ֶY)o�Z� �Ԙ�'VnbĮW� �M�d�Jؠ�ʾ:FʢȆ�2tggPRiG�k$U59dna�8A�+�7�W�9��|PYe��!(MoJ��z7�-K<�O�A��鸡w" ��)��"���:��Y'|y=�H�I`ȏ�O� ���C��T���!�<
�o�7��)'��/�]�����ܞ��O��(����G��F�
bܽ3h��{	�t����Y� �0C�������{�D@6&G���_NaA��2�:��"�;�/�A^�\��[� ��s�p�_5����؍U���k�.���dg�	��d�Y}N�/�<�m|߆�4�*j��jW�o�K��p����<�����2ߤ��Z����ٛ��4��x.\�k�t��]b�}"IbՌ�M�r���b���Mg�>���\�a�3^�D�/��<��\Es:lNjaK�"�w��hp�A��1*�x��ۥ�ã�ַ��}N�h����5�Mxqξ�;�R9��e�e��d4,���B205D>؜�M�a�ӹ����Uv��5���4pC_��=���;��q�6�=[g̜$\W���� �����
	����u�6+K���H2�l	�23�B]�����|�L#gy�Ʒ�X
��b�er+3�É���H����j�&�(�)�KH�q ��[@�怙ܾt�l=%�lc�c���X_)6�����X�tgD	;�-����kMk� :���BDO����@y�@�	��_�&O���~�7�S�����xC5����¨|�o���
l*�o��w�o�����6mh�_!/3Bq�w_�q�\m�bf�[�l�\�È��=�w�뤌�&�l� �����pw�iՏ
/º��v[} �Ů�8�Q��X8�@8$�h=qw����.Zf7��1��$_�%��$9�N	��j$B�Z6��^�������� Z�l��8�˄깯c���NP���J��_O1Q����k�Ч�L�CW��?Kgr��&Ó��A�l��	����h�u��ɩ�u0 N�\;�~��J����5k�w��EP�� -?T�~�8&��X����w#�6�h��۫���L5�f'%�����7�2BJ����}~�%E��)��_n~�j��Z�$	��Q|����Gq�&���̃����:��zIXO����*��ή���&=��Bf;���37І3���P֛_ :6�;ᬇI��5v�|Z���ЭM ���^��G�4ۙ�M,���}�<ϴQW�C��H� =z�7���ؿ��r�y���F�F�^�z���J)p�%	�ME^��{�ay�������Eq�'du�D�ڙ����j���!�釲�F�� 4}����wni~n�l�٭�%�oO�Q/:Suyb�:���_ǘ���	0�>��wY,tYU��0�GQd�0�g�����
�&����J�EABT�$%�A����Α�AE@I���k���" Lr��n��������\�5�s�s�s?�s?��<ȣ�);@ůӯ4I�R����k��=��{����J�H5�՗(�<M�q�w8e=��^��~h3d��Q4��'Ȏ�/��0���~��{a����l��� �����I����������q�~qj�((�B�N���)eP՘s/���l�6��)ы�3�nt��T���T����t7��A9kgz�9�ګǟN�v����GsxE���kmЙ�!h�s�q�PsC�ܡM�D��feF؉��l}�5�X,��5+��x׃I��Z�Y�J>qbKv�C����T���K�X3���ː�3�1��'�Z�[�;�{en�ݫ����9~�5E�ij��M�t!.D
��i�tJ�|v�j�ż@�!��Z5G�1�,ļ�� ���{K/Y�����y9�ߚ��ܧ~k�Na��u�
����IA�O���tjLR}jV-4e���}�$%��t�^sXSq��4(������)���bq뒑��~�S6s�M�K��u#\�*�-����I�ⴱh5���P�d���܄�|���A+������R�ue�#����:l�r���J�UO|P����t;^��/n���x�c0���Z5q�ո]6��gI4d������9A��1n�߸�?Nţߩi��� l^0���+�A\aB�LCp�5���M�uE�7]�?�Q?|��g�ib��K�ި��h���^e�*ذ:�R��dC4�ks����
��sWy'�����k*O����3ˋ{b�V�9?��k��y��R��ˊ"_F������e��F������ȢY��Q�W[h_����ox���KTZ�-� �ma��[��ߜ����iT��:9m����I(���D)�y��p�'�1�	c����][�|�S��}����ϟ�F��<�T޳��4��G\�;� �4+�3��TСP���tU�|R2����������iF�&�4k8�_rͰ}�T��n��0l����O�Mo8��҄Y����%�^��aX��a���W��BE;���.��a�ְ4�[��ȆF�XX�m���K��e�8����������Y�\/v�(m�kd��#�~%�']P���m_��GtS=�:�qP��x�
譟հ�(i��m�1W�}�Ѭg@Ȫ�{pO!�=�L8��,�N� �2I�#W�ܚ�I	��`C��� O|!y����G�i��t�XHL��.f	A>}����{"Zw$��O�j�����;�D||���؏�!s�L7�,C�L�6�P�
���_�������gse3�@`?�i�>q{ǹ�S���L�h�Q
��� �km�QM�V��AsZ�)ҍx6_��x�/�Ș�G��Z �!h;�2�q~6����~CQ�O��$�16�?�[?�F��@߰�N�@q�|ȴ�a���@���F�*U�FU[��%݄ "j��*Qp���mΣru��
�l����Y��}�旾��
~����N�8Z| ��X���GN\�����L�!��=1�n}�y��A�X��CIS�"vcJ[���T]�R:����O$��U�7[EeX�s�( 6�ӅH����g0���"L�g�����ѳ��pjn|���8S���}��N�\F�V�,~~"v65*�^غ�u,��>tKo4[�RA�eB�C�N��JJ�?�0��(E�D�E�s��6�\��|M:!8�v��g�H7�τf��PD���L���y'hF{nm�<�b��7���M�F*�CO-dP;F�h4��'�R�¶Kv�1��������
��^/�K{��~dkb�6�0���X2�����P��<�O�@�`��U ��8��J5�,Vy6�������X�mܔ}GT��D��5i������@VlQH�H�n&�������)�?��c?�V=m��}�ɾ8��A�Y��I<�io������Q���|��8ä��{?�:u�0h��_%V�)����?:��ج׭�>��9l�BG_����V��]�p�C,m<6�r
�sz���i����`�O[�����c��/���H=88�f}O���

歚���;��	bn�QD�5��%�l��_N�����`�C��l�ƒ��e��?S�6wGr�	�hF�����k�C6A�x�h<�xv6~8ee��d����2져����w���+���鎖��ke^Oye�BQh���M�J���ky/�K�͍kS斉%G�ڊ�N�dp��F�����m?� �}f�[`{��Q�Q��2���!|O���hRc/v���ܹXS�&�'���~��^�[Ŝ����~&gg0�n\���Ay؅	 ��H���'cD��^������>Q�
�?e��M�Vg�4��]� X���xTj��9Y��`JDө��l��q�<R��'y��G�	%R��T�?.���]ށ'~oB7���_X��'�ŝ��~�	�p�����L����=N���0q��TUUGY�^�
}hr��Y��Jb�s-5btlynܵ.�YW��%E���&�:�������`85/9�`!�g�;�^]�2�!k4Y��-��PN`��e�rk�s�L+}Ҭ���]sJEwaV�����l `��G������������q.��4�3�Q?���>�6��l��di��\Ɲ�Df��F{��:�b��yu��܂N)o�a�g�m������7��5o�����jy{�� v{[ޣ?�~�z���ǘ2�e�?������PZj���N6!�S�H������[�N��V�|�'�8u����_D=���7�r<��M���儎EX�_��� ����ω<m�m3ˎ���L� ����d��N��'�d�`c�=1��L7 <=��(U$����h��_��jB�C.Z�Zu*��<�pT4Q�:�hB	eS�0E���E�#afIA$5;	Al�hS=����A�@_���X9�<ĄY�[�h�(B��Ukܻ~}e��B?�VNJN�9A��
+�mLtN��Ʀ8�xƧb��a>��S����2SPWu��U&i�4!�_YE��#�J�J������g�aN��]��^�le	�!�1.����][������P�k�C��L�@��������rӘUy&����<Ys���P��B�XZB|��7mxa-����:�#��o���O�@�������`ޖv��C�E̰>��΢�=����'oO:�,iu>0!H�-ּ��\xDo�'��`�:���Y�`7����Vs�Rޒm�G���D�+����摄������s��򓤺��a��Z�qN��{�R���l��nR?��0S�j�k��tz�gT�J��BH�'���oǧ����4{��U&�70E�ƫYv��Tf��a�h��~w���'Ɠ��T9T{��&OM��3�bi�[=�w���Y�.�\����� �u�ynZ7Ρ���1Er��&3B�/ڿk9�%e�G�!M�'7����#��<Ծ3za���ة�� !�ka���ʓ��##�i���{���-�����4���L�㔛����;��cv߹Slэ&r � �o@�B7J����vyG���S���k��7w<W8�<������/<�cai�|&����9�ɝ@�N� �p�]�)������zݽ�E����)����8Ό�h��v�R���Z0�p�v�;�V3�,��y�R��1���[�߿����p�j���Cb\�C�΋mt�!q���
��N�Z�^����녒� 0a�U�G&��?�'@Na��}Ί��^�uܤo����_ܸ1;Y鋓�fX�����s>n�����X�Fc��m�7�t�R���R�4�rw5��C��ř�Kz�^�!�Ĺ݄�H��G�]5b�%[��1��g�?�pl,>)&6�ߢWC4�Kؿ3��+�EnG�{��N}�����o���k�����8Ojt^i۬	?\�H�|�-̍@M���u^���k�j;��j��P�q�h�A0���|S*m��p;��uC�$��3gS ��e�Y+-Q`��C%&=�X��x�
4�+n�`�ώ7������&BE���T����&� ���'��#e$Wz���0�V��J�FI�(�Ѳ��/��Z��D�u���_^��;<�e-��*_he)�^�YE��S��^U�����ʈR�&��vxӣ�Ns<Ȯ��+���n���JT���y6���k��<N݆�=fK_���N�#���Us���r7��@#���ɥԝJ�_�N���~	xQ`�
���ˍ�oY�R��Qp�q��~v���Mf���Ѧr�>Bd�zCt�Y��Bݦg�~�0��~��R]6�E��,uX�M�b���aG�jΉ�p㗼��o���[�u~�%:�
�Y�%4~���sLt��C��Fݣ�fC M�<����ӣpǶ@ў&W�?��^ۚ�rJ������}�61t��4��{�&��XKvm�����
����F�%5�[m�~�M6���AN/�Ƴ�8\��&u���^o�\��;c���5���D
۞���k�8����f��3�=VK/|F��EX7T	����U;��|1�b>޸�i��yk{@��6�(>7q^@�.S.8�������!���~���I��^tn<���{�p����w	$���e��2�Z��D��!I���3^�F�2��3��@:C����u#��˞[��C�0��$�_UA1�i�_ZbD�AUǧs���KM3�������j�}]�ܖ���=�憩{E���?���7�����_i?��Q��ӉM����{V�q@���C�mo/���/'�D��˸ ��$Z�?����'/�3�"�`��e��J����=^����?3|jD~A&�����<�d	�y�ƻkO_n^�)���g�e�=N
!`%���k� �a�醲{QY���� �� �����ѩ�,��W!�cm������#Q�NJ��Y���O7�l��m����l������c�gk7O|l��n�ے(���~M`����A�������W��G	��]~#I�r\B�ˬ�NH�qω��5�Կ)8N�T�[C	��+����H_���M�W��Uf�Ӯ�^ؚ��\lE<m���'dGܹ��v��w�w��<� '�#���bƗ��ѠNx}ه��R�=K��jD[tnz�o�Mt!l��%m(KC�b�JH��Jl�҆6/N�EF�&�����Dݞ�[�u��s�1rV�x���̿y�sݥc��� 30�Lm*�{��2�h]]��.�$�)uS>k��y��١�(��`K'���H���}�?���z�[?�m�o������ZT�<��8Ȕ�a%�5"I���O'�c=_:��U�|A��:B۰ǂo��JV��U��ޅ8'-W��|��+�m.���Vege2Uo��X��*�v	������7�|�v19NMSX�}�ST/Y.����9��<�hIY�^W ����.���t�S"S)�b��jq&l�#b3��woHl��z�	%e����{պ�lD �K�����?�`�i���&Kg�8�Ha��*r�%7��F~��N
�m(�����Mǆ���߽2駟;���[�o`�-��hM��ש�a�Afv/[Ak`/$_I����ۅ�o�s�w,���Sl��@��?[�;�8�@l���8D��z ބ�i�q#����F�w6�[ҺF�Y�,�Q�������:&�;Uc���|�@�7��R�{o{���@�G�O�wV/y*1���[N���3[�L8�sc;��D=s�z�+1���]�;��9�2�,D #R���G=+�.C����B��~B�GY0=P,lbj�[(�oeB��6�yؾ�4mrЁ���5S�]JJ�����MV�V�a��A�b���,����1!��j��m��$�%�����s>^.�V��KJmv�&����N/>��4���Mt���Ȟ�|�K��������ty1�4��Z��GA����֗�wq�O�|w��x޽'w^�x�w����s5�t�����m˛p�5ѣ*����~*��2G��<̧�������hKy���|��<�Y�K�X��dS�a�z�X�N1��Zyp�ԒЀ���
�9�k�����&�ּ�?���3�����ŕ�z��M��H��C�o��➮Ϊ3SP�㴊��_��J�W�f���DQs����F���1Ð��;�Oɺn��#�U~g絭�=m�y.�W���袤c&_v`SFS1�d��gjw�D�H2�"��i�AbFh
(�sn�t�9r�FQ�x"/�1�
⨽/s�5����<
Y� �ذ����R��8����'��5e�qX���d�����T@~[�pi{���)���Y0MoJ�,�9��bB���v���8Z�=#,��A��H �n��6Z�BM]�<�r"�K�z�>�"��ӹ�^g,ؑ�7�6~BBI3<���G{=��ۛ��X������/@����X�RjF�6�r�����C���V���R�g;q�օ1����aR�dԇR'u���G�D��p5���|�V=�O��lސM�U谐���f�0� 43мU��We�^]9��m�����L/�Wﾑ�w��&`�����6���I�Zw�������D󖰒��D1[�~y�N�Z�N�w�g�IVi�O��D����J+�/��,7_��x�2��}�o꺥�|�_H(�1_58)�*3Ū^H'��6�?�+�Ϡy�8�ã���:�jn���v����V���3��}X��ՈT�$2�0��?,�����iw����
��pBN٩Q��=bi��X�6�ґ�'w�EFa�3�ub�V�JJ�������_S�Q8���x��4�*V{ �����`�F����i9�y�����2
����'g��U���T�&6?"�;->G���Cr%��)C����TPj&j�*[%�b�\��[�|y�#IC8�LK�Aރì��j�Mo�&�8�� K΂W�HYc�ü�J�M�8�ݓO�"p�n���r�v~A�'�/����tK����["`�G�	�6Rr�-h�:|@r���!��R˸�G!����g��@��h���mB��ĒҤ2(�H'�dl�R20F�^OCi����u�c�5E�a�&=�<�Kwft.�"�z��>�9L�Y@-�(1���G�����HPXص�v �*�O0�tӛh(��n�R����H�E������e,�DjG�5���ɧ�*d�#�i�_%�5$�o�2����I(�����A˦GkMOL_6�
%���K�7M+?A�<բ{⊟)!"5qIC���p���ZuR�^�<ԄrϦ��n��L�~��%��d��(������&%G�P�_�:�~���aؠ;��kI%#zx0�ˣ�����2����\��1�F*z�^C�n��X�DTU��td���*P��Q#�_�9�(ri�����l�z¤�]W�#���4Y>B��x�T�����s�W��b���y���EV$�}`�Xz��-M'xE8W!�3�5䮔��y�T�=�y����x�	b;jݥh��AtOJ�bƻt�'z�|�A)X9=�� }�3N-�"B2�/�u��J5��`���q��(�v�4��"����枱6w@>�0��@�X}���E�W�ϭ����*�R��t�X���N�\�;�
�Iz�=[�L׺��X���U�:Hbjۜ�l�"�l�?"���o/@g��Ss�3��*d�,症�Eۂ�D��sg��U ƚ4ȡ/+:�,μ�ݦ� -bT�O}N�u�xU\�X�M�d�M�GU-�j��w�_:�|��"�>��L��$V�31l=����,�fb�ߡ�*����� ��M�}��x������~�{b�f�c�~�����f����҂X��Q]o��
)��	��Y{��3�M�jY4|]QwO�{��R���8�̲tV�����zh�;��v�1��]��V܊��0�����?��-׉����#>]�_l<z�"�0}���h'�9�n��ϐ�#1	ɞ+��<��V4N⽍a���UQ�tG�(���H�הZ�6��+���yy(s�@�J����SgޫN\�.��*<�T 5�|&h���G�cJ��-��k[O>"�jݏ��z�y�kS��U����!;��O;1�!�o,��.�wY�Qu1Op���Pֿ|y|��ݘ��^���j��s��g(Q�z�2�������;a�LH�E��=[�5�x�4y	uJ0OT}�b�p���gM3�6�vU�.��q^�w1;pnKײ����V�Q�:����& lރo \Z���C��������p���ZuP�8�D�7�
o`�]PE��ٝf�s�n���v�+N�!6�)�Ey�6�9ž�[�Tu(e﬎�Q0/�-r��2�����]}fn�!�5��� ˟/�x/�������?k��"yH�^���uZ*P6�����Q-Opm��xZ��A^rF��U'��� ڮ3zK��/ͬȝk]*�g�D3
���\��Vtھ��Ɲ$�"5D�Z_DH��I���HH�~.mr;��ߛ�V��P�����3�n��j��$KN\��}{ f^ 
Ǯ>y����p#U1���0� ��t��L��N�*��_���מ2���뵻�S��v]��QC�"�\G9̞���V���,����k7 \�8��H��A��Tj�<��xL��X�έK�y%�t�)?/Ya�d'y�xX�B�ާ �CѴ�+�T��R�2����T�����"���p�eA/Y<#t�����!ٴJ���d�r7�_��k�
�P ���]*XlS����3b38)���p�B�J�5ĢR�a�+�;,�n�X'=����7<���z��PGI��9��_l�Z�p�z�XL	TTn2���uQ}���Z$\�Uw�C��a��PXwT���q�V;��͛��	bQ¹�$q�VHpV��~�K�c�喅;�wὪ�x+#�y������w��z�r�qC�I��n�~��ۺF�Aޢ}��g�q,�F�nIy��\�� �_�|�sn4�R���S��Nq1�ub��1ǽ�s+�W&y�Ǭ#��ɣ�v�'��-)Q,R�L�����Ǧ�_xfv�� a�Y9�������۾'�R���`�/�%��b{�"�#�v��m(�^��$�6fa�������x�-0��F��G��/�c�ʪJ9�1�P�8��$>(��[v�B�Zi��c}^��z�X�Z~X�J���J䍞�=���<ݞ8�:����g����y�ɜS�bõ���%ou��*�p���r�jy�#�XQ�{1�գ��J�������nCz+�de��қR��lx}�a�X9�yu��9J�m�i�d��}��y�1�g� ��b�e.�` �l�y��S/��pPy�g�h�n��՗�skL����R��GZ��	�9J���N<����}������f������N�"�D�6���/h}��
��
)ٴxZ�W�w_Y�:�ĚdE�.���~^$�|ʰ�������ݞ_Փ��.8�gѳ�Yi/�E�W��`��E2lS�a�$�[�w�[-{�����6Jm��ᇳa#�
����ڳ����Kߠ�X�R��l����e�ɣ9d!g�����a��cǐ��"CL{&����e� b&�@�*�������B���q���ɾ��P�.𚊑v��РQ�+�$��T�Ğ��O�����.OܨD��M���s����|)������@ō�@֡�b(=�*=���8�\�Vq=�0l5�s�9�}��K͎T�
ѵ�§уD�:I*�K�.�jJ5sЅ��'%�|�a�,u�{mM��C�����[8Z��2KZ]7@�@`����v��;j��\aq+�IEO8�^��K]��Smឈ���O�&s�vru�e�������sEd�使��	?�R^]=���c/�O�fř��`�*EA:\V_���^�6��5)&o����Y�*ϋ4�[S����fI�L�_��8���$چ��m���d�:-	;y9�L��J�Q�OR���y$ߞ���U��~W{lpT�f}�\tyB��k(�z\��S ���w&^˷N�ک�-oz��$J?+��ۇN��H�%K�:I��1�W/��4���NOg܅U[�o����E���t���.v+�>�6�����*����V�P8�$��և33�itH:<���8Ή��YB- ��i��.rr��R�+��WkE��r�VZ?�c+�	^s���p�͜g�hk2��AڟnvuM�C5^7���.$�4_�B��k��$���`b����*-n���?W�Oݥ�wr�{��u�w��;�m\ҝɜq	��z�w.ʹܘ_�;L�>��`����{�&���aK�B�ӛmeK����I]e��Ip��aE��n��˚���\�]T���]��������S�@s�B�#�R�{���oh�Se�2uۀ'U�+1����s�rf	����A�8K�|(�"��ñ:��c�'6i�� �Y�c$1�<�IѾ���A˄�uR���w���]���l��1�[�9R')t���$h[D~��+W���W��0ʰ\�@6�cVw���6��a��x�zi���<�.�ˆ",��.��V�,�H��� ��9��!j�ލ�?_\�#�7e�b�i��Q��$�R��U��2HS!{+�
�L��[I��{8�@�\�?���_�x�����O6<����Ry�kY����9�S��ÛϜ
�ֶ�ȫ����N��ep���S�������eG�v�!Sj�a��=���Q��D]~(����ҽ�}��-T(��E�9�ѰdSP����X�7�ҏar_ku�k0��O߲�&-�.�)s|r�kp��,9��A�=���ӥ����rK�[ޠ*N�l���|�Pm���C����})
�YG��c��]T	OHS��6ڜ�n���d�ޞ��3%T'_�i�|��2���1�.�mF��d"K��h"�����L���yM�R
k�+8���s��sf��HI�Y�|�t������֜"4
sƺZIz�MR��߱N�����~�H�[^:�;?����>u#r�2�Cs�����4�DÄkuir7��!m£���ѹ�:�L�K�{b��0�Ș�߶��*�ؗ|ھ�&�-���S���W�I�Ê��'�v�w|S�"�MD&�����c�*�>O� ���%b���2�
Y��V��Ƅ}�4����yֵ(����.�����ko��g<D$
�z�SV�h[��x;�<�"V>�ȧk
�p�W�N}ڀcT��&l������7_m�ª����.o���d��B]���\o�*ſ+E��a*���D��P�ž@1�F�(&M!5́rk�_��ћ�	�0{�1.�L,�?�R)�[��^�% ���)Nx��Y�p��p�\���x�*t�ħx|�Kǯ�?"�~EG�ljO����j=*���;X�|�_3J$J��佔�	�Z�,��h%���+��Y�]��.Z��uA�I��˂���6Ź�k��8@%ZG��M�C�C�70*m�ح�`�b��ש�k@�L+���Z��A0s?X�?F%'�b�/yM��'���3Ƽ�Pgp|�c�-�f��b������X��N=mw|�BVծU�GH�1>����GY��!�?��%�������������H�hHn\iY\D���<�_X^�[?���l}��b<�?�ͿBՑօkl�`+k˻���٥��-�!4p����,.\+}kغ�����ϸ�)�z�Q�+�2��送�{~�?�I�D�mn�wV��If����݆8r�+��7c�B�B�dp %(Ͷ*�3��`Г>.�A$=�Kx�إb�Я�aG]V.�cSwVU��X����4�qFT& +��'9� ��/�.t��%B�����;�|�V�3Y\f|�y����'M��7M��(�}���Ol�e��effa�~��}Q>_�������l齃U㭯E/��a�#����������۩0˞�յ��r%�\jO�� K�l�J����M�Â���I�hvD�PHVoZ�� �
#�qym�%�3����A뗬�3�u--�R �8���,�ߚ���A7,b�pa��As�O4�C�	f������(\��k���-�2�?g-�:s�JHIy�c#�=��XL�ed��q��p�K��q�<�vՆ��O�W�����L�U(Ye�9A��
�]����e`�\c�Lfk��&��/�7C�b���Ў���ݯ*�~�w��ե��Nr.�sYcqZZ
wc#aU�7�����S�ږ��{#|��,̊���䕉Dĉ���K��O�n)��/}*��IL��+�c�ǔ�~<�3���>e�-�ǈ�z�|?	�y��*���н}u�)H�4�(�z򈂁�����{�'
߁������e�����a֏g��������Z� �;��vĨ���*�^T��������!�?�Ζ:)����>��������<���h�<�I���$� �|�t��̪���>Y�~��]��u�ŃiZ��H���������>��,�N��F�=�G*l��1t4�����5���nW-#q��~uYlv��9���J����|N���Ҝ�['�d�퍶v��g��Z9��΍��s�FHV��B�T.t��ΐm˔.�4SJ;�r��g�K{v���]�ۥ�}�I����U�mS�W��ߞ���9d�ث��a<����>zy'K�g2�X����]����q�U�}B���2	S!�)�#ϵ�A��v�8i5K�%�m}zu�	�s֢�q���qI�Ԍ��B�?�i���'�;�t�~[�OLstYzUfK��V�a|�B���In�؈��A4�����[�?�<��,}��d�s�H-�)��'�!�@	���럚\LF6�F9�=�h9���5��V���$(���J��k�2X�����v�6Kxt�D4�<��n}�O怳����&Y��>W�T�L[Ssdb"��ނ%%���.���~�X�����v�ڈ"���#�IEcr����9<��i�v'��D�%�ջ��y��b�ㅏ�>*`*{��Ϊ�t��5�,v�+dWe��^��U4��G��.]����J�A��0�;C͕���������L���Z�';�W6��Y{�o��U�[u�k�$:L��O�})n@v��?�=*�;ݗbYY㦸!-�Ӕ����!����*���7�̑��p�X�*�6��T�u�7{�}�9���Zǯ���������[��݅P؈��B	.�D�ΐ������9���d4
�N� ��G�v�c�����`�+K|g�@!�>��*[R�0M�zDI�7|�K��t��RJ��$z�K������~c���K��A�ܩf&���K�Sa����u�'�3ś��K�W�|����d�AY۱�RJ���(uC+ nA��������\g��k����/y����OgP|W6{���_�M�ۈ)w�x��&8)�L2�DX;��#j��O6���Z��/� ��2N8��*?��\����$�PJ�k��̢$��a��+��)	�k�U�����q+rv����驏��Z��uk�i0��u��pRT1G5�xI7�*��Q�_�'S]�#ʿ+^|L%���l]�����e�?y�C��ӽ���5Uꪴ+���K3|��#J����=!�����H.eb�k`6/`�M5&m"`pF�����,G�ɕ�Wk��3B9��sɖV���1�>w~�jVD5�) g�Ř����B��!�q	������l�o ��^������M�Ð�4nE/DoZ9�Ĵt~��ۥI�-J���k~�����N�{���ى_�[�ro��G_����b�{�������L�j(A�4�nr\�.�=࢓�ž{��.d�_�tkbFΤ�B���N�Ї��,+��M���+J�5���x��AƊU�B���w�o�9�>C�Ml�>M�(��|��+<:�ùP�7��ٸ��YBe�+D�?������sʾf��M�!�Vc�z�#m�B�h *ע��ɳ���?��ϖ�Ò¥[:��a;��a5ҖCL_�S�~�_�=�#�Ǐ-XN�W���Q��.\�;�����m��]�����oKw=v��N�=�e�MU���z2����ݺ����\����Ý���d�fL���d675��Լ���fV���DL��2�\/�:�%�=i�����=1��4�3F-�j�7�L�L�`:w��}�L~y����ɺ�nr����t[�_� -�l�	�u~���sgi��h�#���5#h�ٲ�u�H��=H�:�o��j���djW�S�^�Қt*yQ��#O�|
�x��ED>|G�A�&����T�I����W0hu�q����7Ơs�9�*�`}b�IM��4���T��-~��|di*��E}��=�\����&�n[�ʛ�\$�oH��Em��f����C=��#Ak!R���Op83�
��x�d=��4��F0�ǻ:�*q��B���o]՝.��%��e_�٭8�����<gw6��>#<8a�>1-/��Y�
�g�
hl��<D�hE:+ �]�Z,<�64z'��"�#A���ݝ��h�c�cH/F��R���<�.�j@h5o�]��*E�I'���.L��?g �16߽�f�����P�\�:�cZ�;�®˒�?=���;�
Rï<ʁ���ϸ��������@����Ē���mb}&������Og���V��ua��	ZL������G��3������xu�e��c��j��6ҁ�!�o�UF���5�Cb������wm�Nܮ�D[KHܡ���
����	�p]�@�2F	�m%�	k�~]�H/�_莗wm�45h�H�ni�f䢊����sQ�3$��\��G6`<�ˁD�����dm�.�����m���2�k��&��6��A��L�.��r�@	M�B�b �<��}R�.���N�;�A�&�_�����V/�L����dI��PU/0��o/��1�7��Nc�m��.�U!	j�=U��H�`'y��r	B�Gh}�ڪ�K\�!j�� $IuC����j���I����dߓJ7t���6	���Z}
�u�5fb�F<㪸�]��k�����XG��w�#F�깚�
M���N����ͨ��A��Ir�6��H�0j�S�;E���!�y�g��:��YY�O��E{es�0�6�j�����̝��[�O����I/n kU��M-w�#ϼ�J�� .+n��?Ҭ����Sy��:
���}�Ժ9���$���?Sx*���~���q%��,W+8$��i��?v�Z�v�k9�Xs�4���}�(�=`����R&�1QN�;��GZ�4x�iA��8�%����O�7��`1�0��t������V5��7�4�P@��l?Ǒ��@�_F��L�+t�t��.�Y��ΛzD�B����i�?�7�ÊJ3܊��K�h���vF�̙&0��d1; �(PV��O�~�kW��Ax_Ѽ��E�����Ȑ���=V
^����+_flO����r�^3�q���Q��]V��n|Vk*m�񲻨BoD����M�ݯ��Ռe��hhh��TEz���N�;�<&�-��Ҟ�����3m�)�
S���D���Y����I.B ۗ���62��4�~�*t��^�i�?�'k�z[y�b�:Ǔ�~F�竡�ݜ~�6Ƽ�pŭ�{NuDn�&gJ���,���|�`ei]xx�a�u��Jd�#�K���G>�و�QRY[�헜�����@���~_z�5��?+l��&��J� 9�1u�	p	B�J��PY����?�S��"�p㭢��l���%��S�AR�;�fw��O6�)W5��ui�O�(�Kp�*����W�׽a�j_}�D|����qv�1	�to*;�1���x��}�ҪY酯�D�D��'����	fUy^�OcD�P\���;��Q@b%�5\���W�:��dR,p�GZ� �x��)�yUr�]7���+���#q���x�[Щ����B2�m�*Hg�֪�l�I�����t��o���cX�Ũ�}.�y<���im{pc�vգ��7�)�:kU�Qث7ɣ����|%;�ؗqK��Omq�
����jZ��#���f��(�8�l}��	��v�2�H�\�=\���ϔ�K=��Ej��W��>��@�*c��"�H��4�XrPJkn���<��-P�N1{ª����N�ۏy�q������Zi���2qtI��}3*rdc��/IɿK����m+o�V����/
����=�%�b��y&��vu�H���Ck�/�	��8���y�e��$H�`!�LK�����W_����NO|�ʴDV�q�&To�!Y��������C&��JN��-��".��Lh���YQ��%��o�!����x�8�V���<4�d�#9Z1+�������Ur�=w�s1�z�un����WG��n�NL�f���;��f�;(I��K9���U�z%m��8���
z5EMc��p�t.sd~�R->1�sGJxOIpo�qn�?2�~���N��/���l�i��l��@}+� y�^BmM�h�z�������H�6�����F�f\�kM1)l�$��G��O\�(�SǶG�K��<�]Y��(��6@br��$�B�����$��.h��ߌC��z4�Ŷn�������1�i���o�m��̪�����5ްo���'�����!"|��8���5`��r��!g�dېdc� ��T����ո(��ϻ�t4���q�Z`�Ы��o�dy�Cא_��L���x�c	���~�T�uX���>�r��4��E@Zb@Z>8t7���I)i���Ai�������~�0p��{]�1��콟��u�{���d�����L���7�����PY�o���S)�;�`Q9�09x&��Y����%�p�ay��Ur?��,͜�3��~Pu&Ǧm�=Q�\po1��5f�I�7��~���ޥ��+gqrݚ���{�%_@�6�n��̪�ܡ�V+AZ+o����X�$\��j����V,/�$��2 &Y���~�保Oy=�h���ߐ5��>�(� �q�Gq�M,,�a�i��{����kZ���H�0�Oee~��r���Im�Ɗ���bl���Y���bB���wU�6��T/�é<*+y�)�H͞����t����3�F�-�?����a�'�2�*��rS��6e���)Q�[��FH�5�~�]B����j�[�u,R����'�2��5�9����y$��ϝ�
]rq�˓SṂ�9 ��~�O�$�������Q�0 ��~�c����A���ΙYY�q#�>��-q�^���:��n��{?̴��6�����60����Sp�������D}I_�>�k8C?^]w���--Tu[t�(�5�˷C3�>��\��@lё�8�$]�縧Ɯ ����@�緩��Y�㒀�r��^�����f��,�w�"m��`ך�gC��C4s��� }��w�u�Ǥ�H��3�<8$"SX���ɑ�yΨ��L�/5CU&Rp�V�q��>�g/*;���}b����=C~��|$��������"��yͻ6�_�q�pok��a��|_��dW�9����>�j~dX�_]H�]����C�v?��z� /�M������ �,J��|����y��HJ���G=�,�`�r����`x�Ȣ�=��Q/v�D:-�����ыgv��/�Y�yg�Jw+����e�������eF�6�bO���m����"�k�]cGݏ|�oҗ���:~U��1�4Q2�6��<�z��>z� �\}{��>�?�/��8��9��{��1�Pp�9h�W�uQ�'���J�{��K5a8���&��Q"Zs��*MTs�Y��9Ւ9:�/�j�٫;���Z�0���	ͩ��@��ُ5�>Kd�3ZG��5���OW�����3Ym�g.�ۖ36`���2-ȏ�l���.j�t������MƓO�'%0���@��zf���Z!�"v��&�0���6�� V�v�mW����^κ�����h�	�������]+�_ӽj���mYAO���nw��M�rF��4�ء���6�Ú��.&[���'P�tnQ=K#�u�S$�Ǵ�a����w|2���N�Z��_�Ӏ@M���`����qn��
�����}y�;sή�F s�l����WSy� �%�m�
�ͼV��I�`x���k�7�[6٢����D=��c�h%.F08�_�H��u�J)/��R�I�'ڝ|�3��Y�\X%��_��d5lp�۸�|c.�z�\|�6u�x���TNjw�l�޾����v�M�	x�|3���dz��I�q쏧�&��Í�B7"��ji
R;�g�
KL%m�U�����a�ө�Ɩ�����)��2ߢ�a�1r�OA���[��65�g��I�zYuK��/`y�0,a��ZO�Eh�H�4��&��`��"�p����oj/&�Voy�1���|���k��;��+�#�Y��6�]?̈rF���㶵.g.�J�sij���[^�k*�0�ӐV=e/�N&W:2�d��(�~���qu��X�XprV$h/�%�s��!�\}nXU�5o����X"/x��`�x_���Ǆ&�_V���I� A֢֮2�ѫ��.�2Qm7��р\b�0"Y��D��N���{��5#��t��N�b�!ѿP�"���r&�H_��~ȧ|�GP9�,��O��o�&�?�Nkz4�U���oVZ��*)T���{�m�T�ٟ,Ud}o1�k_ ��E~��t%{��1�W����5.�����5ܓA���O�u�Ň�[5�Ø���-�Z�Dy����GA���s#�D���#!%���}Z`��[���STs���3�]AX�M]"�=�"�*y���A��	r�'!*���x����6ɬ����ٽ�~Aĸ#xr�d�u��5 ���i[�������!�t�E�%�!�n������������\,�-P���<_�
?[`3d�r�J��2bm$ 2\�r#�:���$ǂ�e9ʉ�+��@�m���Խ�ؑoG4>+�f�05��xˎ���o���{0\s��\��[U�x�*��i�b�D�Z4t�i	<��KLٶ't��zY%"4Qs�z���Q�k
_��n����]�����P;Ə���$���ik���-���2'S�-���!��kG�m+���9px
њ��%�(I�6���[���	.��k��sfzJ|U�a'�4i���Qa PV��	:�4�A�Ƭ�l
�y6��8��1���F�R"����e���Q�5�"RoR	-�g�ʤwdf|�I9`Z��eԳ=�@�Hc�Y��_�U����(m�5$�I��Z~����\}�y+�����Ȕ�o���,mL+$�0�a�R?�\��zhTِ��n�R��p��0�͙�M��$�S��.tJ��A���d�1S��O��;�}��s���軐��"B!m�
l����gR���Q���^g����ϔ�3=��sy�k�#�y �r�]��w/8�������	�2�l>l0fi�#4�~yN���7f9�QҨ���A��f��`e�	�ԛ��p�삢�\F�=� j�"ݟ�_��WG��>g�T���#M���|�^�Msᙒo�$.��c�������j���O�g-<^�j"��S���~�G��B𱯣G�א��N�G!����\;����>��7�ג�;ݸW,�%�>a�*���b͠�vfȼ����ݶ*��-V�/x���]�a�'h��f�M�d�6b�RA�3��az<�r3'��\7�7q1��ѽ�ԡ��.����5uٻ`�	���*yc�芚�2�)�%�G 
ٶ��5+�"��a�޺6���{�Ý�#�#DQ�98�E�%���%���C��*v�3�"��:"�T�j��eG���) 3}]�c�Z�M�������%���Xa���0�G'-Ӟ���8Ѩ��8:!�ν�eF��f�}%ߜ���QA������}A*�8*̂��;�*�h9�5� �
*�bv� �Ɣ������79���F#����Mw������g-Ж��]c���7' �x�l��D������j��'/�N�Zv�a�K���A�Ҙ���>$Ӽ�����w	�54�e���%�'�I�\y���)�Rq�ಣ&H?+>d�%�h����(�u���VV�8>9hF�f��DAEncv?�@g�]��I���غĤ�ʨjTfG4��hf�w(����wC$��CÂ=�5)dY;{�q�U�Wg>6��Y%zc�]���5)�BP�"@tߜzْ�yFig���Р��O.�d�"�h��ؒ �> �i�
LչMs�Y�(���|.�Uw�����ϵ@F\�w����-��$5�=.\4./C��ҳ���7�V�d'!�[�yV��2�H�L��"C3���Ȏ��j��9��&���I��#� �qAe�ַv:�6&vL�YH|æb)A�La�KX�^v�����i�6�)�ތ��5�o����]����^��AUlF4Ź�O���+wփ�h��?����h���C3��֞���d�j���˽����f��TKO''ƵQ�М�Ώ��ϙ�<EFC�`��|X�����2��}�]A���2�6�����ތ�Z�#�ӑA��~c|�O�"�x��pK7a��*��3Ws��N�.��@��4��4p򩋩����<q��k�����"�_tW�0��t>t˖�����FQ���·�6̙����M��d����~���:�K� �W+�tr���Y�����5U�|��N��
��`�����'�'W��:� H%ٛ�ڰ�τ�Q�������>7f4��'���_���$Ŷ�&5��a��@S�����s��`�\�+����A,��^��L�c�
F������T�S˛�:{8��׷�^��^�3`�`��B;��8iQ�Nt��x�P�<m����vaQvb�@�ug�:�|d�>&����Q�A�� }7�-�J8C�:��5�+�����yC�%��;A�X�e����͊L�I�ݐ@�#�J+�
1x�S˛��`�\�@q�J�p���Il*$��ypV���	����S�yv1�b��a��s���gi�+*���1��Ig�����u��@P�������o�J�/���[�t�p;oK��1�|'Ųa�������>��2�+S5�{DK=��J_��k*��mqfg�ֈ���X'N��&�d'��S2����/Yq�s=�3�S^�;-!ݓ7鬠of� �D�/�j���J�9rf�}O�:�T۔��	g�3�O���T7��V�b�.�1�$�-Zg|ܝ���CM�x�u�B�$VW}��3��oLF[hzR��UVk~�Ѹ�I^�ɜs,��B���8�8��������D�Yx�1����SK�G���T���k�T=4���s�ܣ.�#�aZs�̆B�,�{�*�E��&=:T'��#�Y�7j���U]����zO��XUH���C���'�����QSǲ�A�Ep!�ْ�J��W1�Suʍ���X�Ɣ\�ap��ze8�Pt2n$
��4!��X�Z��H��޸�>s�������U<�-����$NNS�+!�G������2����"���w�<zQg8t��{�;(�b�=WDf��U8d�ꐖ�kd�����؃������p�]M��J�V�E ������Ȳ�<���'>�zXT�.�����HCu�xw1��fd��$�l9]ubU߀ut��Y9��w��V��SXXM7���oD�DU-�Z���"�s��[��� �(.�Z	/�7r5U��k^�9��H���Y��c��a�������ND:}X�>�ցw >�+�����p��ⶅ���@�a1Ɩ� 6+��׌� ��5�i[��a���&Ph���t��zh߂��E��D���xz|�g�tTq�/��������s̚QR�P��ԅ}G�#��АA�T��p$i�p^>��WM7G�=l�.�-kN�lq�z;G7i-~�m��~k~>���!I=�ku�eg�	yb������|>��l������5��	��&�ɱ̱��oO���Aό38k��g�$9��n��P3v�����l��s�mQ����ګA�`���۩7� �N��̶x�:s�쐵~���ޜ0f��_b9�9�K� �
�a\��V��#��)� ۂO�R�\�A�1��T���i�{~,�v:;��#U�O�_������-�~}WQ.�&G����O�m��D�I-��I�Zsmv�-�����Ί���{��!.�yx�\
��i�[Eo/l�/]�.6���G��?�A�s}�ڥ5̽�]�T<t��h��7�0d�f�*ɰ4hµ�fҗ��ԡع��S�d-d
V��Uἂ���o�a=�RF#�P���L�<Kn�`�V���~��.eΓ��u��۲H$�~�)&7�x}��:/�>0J7��uaB� ���S��4 �|VFDjp`�D��e��0]e8*�������1�{d�����H�\��ͭ긁{~J�������lP�0e�,����D�Kd�"�-ʃ���:7g��X_7y<�1��3��SD[2��"�|�7$�o���܉0^��ڼ�s��={�L�@���7r�j�έ������U���9�����} i�Ah�&+l5���G��p�@wg�f�Il�Њ�ڢ��+E�9EoS�ݪT�K
ª?�MvQ7'�}��@y���Ug2��6^�A�8�����rP��k��饓g['�����"ֵ��Qg�r���]c6���a��.k�|�x��U�#>U�Ǜgoc�_79Q��}}�ˋ����yNr�!m�2��TNjց|W4��ޢcr��
� <"<[��.�Ng'��o��I'|*�����O$���|K\���NQ\jԥվ�#;Ra���[r���y���m#vK��d���9��']�_%<:�&m�s�>h$¯���>�.W�*+dEںy�r���*,�Ճ��hL]M
�GL�<Ts�<�_2�̊����Φ�cl��y��k�#g����V%'Dc�Q�^n{��$r�K#�`Ҽ�[�'V��	v�J���������.2?�G m�W�k���w:ZH�G����]�����(�+\��Yf�x��p>��X|�8]�ap�5? ���)Mv(�`:t�����nB�j���\�֒�[�w9�M��N�q�,j���eE��F!A Ryt��8�e���?��{L�Ԗ��=��Ƨ.g\6F]挓a�c�r	#�QT�pXP�.�QT��f��A���G>WMW��G&�&�kSr�"��J_L�����@�84��S��"�)b�0��y��{O�([ޡj.y����_��`��9s��S�D���I۔�Ծ�r.f��l_�xWA�g�R.
�۹��,�)@�@�U#<���N,��U9�zzl�"MnϥuQQ�Q�L����{�w�}�>�A��l*�rW�>��e/H�z_7�0�"aL�؟�<��������c`pe��b(j�����h�"��3̜u��V������٭�t(L"���e���p_NR���Y�y����� l�Cm����=_����m�0�]=�9�w4�d5`��z${�w��r�|����>��=M=E�WHQ��ɵ3���k�b���*�>�!h�E��s����CT�U�����A`�w3��L��X굜i���A:Yd'M*��"����dU��*/�j��}��Y�XLV0,�i/�����$[��݋��#���׾5v�L�w��~U����띢^���V� ���FV�:^��D4���P���mR&a�I���y��1�r���K�~�l��.<�25*���7��3�r��8����)�dq�XN�(Ԟk>R��M.ڳ�MM`c�o͂�F��	��u9�z����*�#jv{)C�]0n���"�����P���ݩl���EG�ݏ;U�i�3b,j�	v$���D�Pu��n1ŠK�2rn��ҵ��-�ˍ\�E0�B��p�B4�5���p��W^ѝ
t�7u#HT
۵L-U[^=K��Θ&HH^�B�z	H��y�|����I+�vj`+���=D�_���u�w&z���|g�0�}� t�|cl�kocӎX�����B�n����G8�D1�DD-���n���D�g?��6/&���E��np7�]�OK�~7���ɎH��&�uJ�i��,��GJ\,�MT�\��M�֋+��r��4N�m�Sv��'93���>�O��kqKZD��_��:"Sp倾D���Z�o�SOS��σURϣPU�P�zg����Յ}��$q��R?d8�;K\�#�?��	dF�`��Q��Q�i�������P^q��' �H���� �����z�:#�~��mw���v��EM�#5�{�[�d1%�b��?h7|�q� \`��R�d|�?�+7��۫5�G�����'��ݓ��O��>��]˻�����X��,=�Z���8��ˋ^�����).�Μ1p���l$v5�H�TQspY�����q��.�@g����QB|9S�m���"�����Z'��暟J+�1�-�Ը7jq���]�t*N���_]�:m(���J^��s��@;��q����#Zm����KZp�6h���s�4�~\>l�ށ��A	�ϻ��0X���IhB�����g�������w����0F�7:-ܝB�h��h�*�6ǉ�vW5ꔊ�/�F�d��I�C^�~�b9�G��%�E���p]�&��Eg����t��Cԛ��vʢNsNЩ&s3�峒� ��� �h�;F�sx\��Eƹ�	3�o�	�u>H��k8�	��{C�ms��9�rB6���M���/��G�W"��$6�V��~��kSѱ'K�o�:6Uc��dy���c�����VH������gI��N!�Y;W�=4+���r�Mp"܈��"���@?�=�����Fxt�?*����S��9 �t���U��n漓#j\�q���f��,�þ3�v��mx�'���P���rv��I��O�*H<"G	vY9b~~4�ymt�C��9�rz���a�Кm���5My�� ��_?�U5����1 �bd+�����D�LOq���� �Bv�4|kI���Z\S���j\��W�D��^����x�r����߱J�_��0.�A��f�إ�C��|�ڀ���W���V�Q�&}g��z�ј��m�-��Ҥ}��oj\�n^F���c��Z.o��[!q�l.�����()<R��[С��ۨ�keU~N��nT�8��αR�����?�na�O/7%�I��\u�PK����W���$��ޗ�_�dMX3Z�t۴I��񻄣���i[�|;����(8���q��a ���f��UKq�Ĕ_�eL{Š׮x��ob�Qq�n,������{�E	
���+�[���`}�+�^���e�#�����2��Ze�D/W!j��K�uA��1�q&����"��vt��Fx��Y�"tj	9�ף�I/����	qf|�|Ĺ]�����l4�ȫj����_A�'zT��`��w.~k����y6��d/�[rv=� ���Um�E0q�x���O�^�˟�_�m�/&� �%��ca>� �񨽲U��\s�ҥ�(�&}�i�0�yI�?]�A�"��q��b��ȳٞ�f�Ffۤ(H�K*N2��,���/N]$�oh%�.>�ݬXLS�J���
�-fZ]U�]�(�ڭ�����5="�X�xΪ�{��g?]nTg�J$\׾.��'��A#|��i��O�![Qշ�	ַPV����j��.B����>�k�:a�̳xC���wK������>�pĘ�%:�a\K�	MY��"���k�[G3dY�:;G&�韖U!`�\iv��O�""��6Y�n��h��1O��A�\.t����P[���P����6R�u]X���W�o�<�HȓJ�ʄ�,��)5����ڪ/M�GK��S�Ӈ�3����t�i\�nݕO�襉���x�i���S�J��K;Z�w���>�.TIܦd�>K�DK)������wG�<ђ@\W��L_hRt�3(��N��3L��z���s���$'�?
�m}�`����N��=�?h����� �����c4nK*���\F�J����^k{�c߼[����P� h1�_������}V�"����^��0�[r��n�%�g���)�o_c�v�{�ȇ����K���S�u^br�{.�ʷ�10����~�+���˭���8�;K�?��=�m��I�H��ß`>J�̼�Sy��>��JoVԶU�?(���B�Ol�� ��v�p5�@Q
:��Z.��,��zow�����XkE�T���	���\뎯�Di\�w*�|�v�=�.���Ĺ�J��~�A�Ït5l���3-�����8�����`�Xi�t
*K�y����).q���Ϊ������f�ɭ"4�'<�
�1���u1R,'Su��X�{ɋ��_�܄��R+r��5��=�ey���ݘ��Dh2zHuӏj�$t��`��[�?�%�K%�j�B]�;^�%��|�[��S�SD_Y��Tږ�+�~)�Qo�1��r�F;��2�9��i?��MO{)�=ޠ.p"�P�M�C|U1ss��íT4�+���6��O��"�)�z�jW�q]��Zi��4;��a��w?
N��V�$�.
�~���o�y&DJ珏n��Fx�M��gc�3��Go?�8����e���\�����Â����˸�����1�M<�l��D'?�4�F*\rT�W0��x��U�B2��6��{w� �����J�~�L7���WR��GL�(O��\��6.8�i*���x�#�]ß�#� ŵй2s�(ƞ��)�W��w�Hj�M��ӗYA�O��F
�φ]l+�>�ryZ\��je]��(�ku��O���*y��ٸ���g�ۮed*$�kR%r���U{�'T��*,�*P	y.���M�y_~%������Y�ɩ42/a��5�W"�����].����$�����E��ZL��^�8l��X戴�� �0o���,��� �T�TՁT��Ʀ�����;gM��I��Q�E�<�uH�]�!��R�ǤSZPf�yv��E�0sɺ�a"�دpt_{Ɩ�rm��6�KVh���u%}ݕEz(��Q
���/|=ƭݪ�B�+O[D-�n��>��6�N��k�o�z{z�Ϗ"�\�_&�L��Ų��g�2��F��}����B���V�2�j�ו'�ڌT�l�U���x����O���*h�r[-Y�l]�~���ɾ=+Q�&<�����i���X~�4� ��i�I'G�M"�m�g�
���0��?�ZZj���^����}|�R��Mc��j�����M�%i������nE+��w�F_$� =��[�\��E)����p�71d����u��?g���i=FY��{cW�[��oFdd�>�.�}/���(�����[y�mÃ��]�$��99Tޣd�+��w��/�7ͅ��<6QKfT^������I��#ȅ��GIl'��^�-�o����C�ru&vN�"CRٱQ��C�����QbM�-Ȳ�<�-^-��׾z��JӉ聢���cq~�~[jƴ=g�QA����D8�'���ٔ��5Q���5��N	)����8�1:L�P�]/xu������Z ���ѿ�_e�m�!<#C(`0��Y�����V#GYt{U�+�+�{\��ێX��(���u��*7~�.D���UX��-\0�]Û'~���k�e@ߛd�rf�/�5�a�"��Y��&xR6:1����&{��X.U��⩐�੏�b��7ow���"y��ʝ���ˮ�D�!�&����=g������d��������kcty>Y�Z�A����ȔT�_rA�%���{�2���B)epk_J��O��qɆ������oW6 �Iq|��t碗�3Hv'���{�z��D���������!�uY5�%�33��o��<8�v��kݵ����i�;̢@r�g[`����x=,S2���Z���nE4�V���:_��G�����BՆ�m/b�F�bJ�R<�כ�P/�υ�&�\#VE9���+�ZE8Ɠ�i]zw2�$9՗4���Xf-��$��~\�^R���4�&�N>47m���D����/6:�_̈"T(��XA:P\T�SeO����%�q���^�-����uo����or�`M��'J���#�%?6�~dS#�cW�}}��ަ��qF�H����!�Πּ`�
s�L�Ujy=�s��F�)�Aru@)��&34�����wOH
�k�AOA�Ӗ��n��4J��Gm4�Š�b��H�����QJ�0�S�*q�ޛ��������Oū�58}�|%����W��~�l�G~�VX��
UᣙOb���ǚ�):�!��y�p���"z�%�V�������Y7e�e�L��adGxB�O����u�M��� ���A֐�q�$����хA	��țj��x�J֣ʊզ94���!y�%��$�G��[�i�(J���i�3�u�]�.�t|DU���c^�Lë��DW��q5Bg�2�挢��j+V����ꋻ39��Rϸ��w��׌y�œ�'�en����Yd�PlV�v�3�5oi����,�MJ���;��0�.�}1��L�4ں��E2I)z<����_�G�Ob��@۷�.��IV�����nsJ��_��)��{�K~О�+j�Ľ������F�8t_aa,0�4���b�lñ^�l/�v�X\Į��Ԛ����Q��U5�x��7�{�59�_�{7�b��CFV�
�8��LX0�*�O��u:)5ꉠц�U��B"oݫ�z��Bo�$MX����zn��u���f]�'3�s��;}��H@���F������ڕ|�&Hp�$j����\:�����@b>{����eBטˤ62�2�
ʎ+�F,`�V���N���k��D�6 �gXY�U�O����ٚcO���H���>�i���g�t������u�l��#�*Ņ�e�B�����FS���%�A�;��u���@�ll��c�Z��3'���8BD!�Ǩȓ[ꃋD@��pW@� D�pwd7��>�`�wp+M����E���vj��>��Z�����30j=u�գM�a{<�ҟ�9R{����K���~�"<b/9ޯ�\%�%'(x���_P���t��b�"��l�0^��z�D�6�z��F��[�m�f7����zdN��J�:�5#���p��9ҥV� �*K�U@�ظ�HQ�1cO7�N��ƛ4�c�HA�l��ۏ����F�.N��ץ��i�?�ɋ���,�M���}�b�XU�D�y�{�7"2D��� ��ᮝ����@j-[5]{�ą��k�GM����Ή��'�6<��~m>$%�~�)IM���%�@
�#�.>1�.o�ˇH��)C�����u������S�+�R�k3!�Q7�4���?���v�M���� ͱ�W��Zi�Zy�#G$̹���_دӕ�7�0����w�<B*s�
r4 �ۼ\qq�/���,:|�oӍ\���)�,�~n-�ܟQ{�;G�Z�����y��&帉����Gq�W!�}{�|�zӛ7�d)i�w�9�~��1|��/��3g�)�!k���C�N�|'|�&��ͅ(3햄M�l�B:l��؄�xѠ�\��$A���<��%|P{�[��4��!Kc�wz�X��P�������Bi��nз�2]������o�~6'��nX��Wܝ��ř^>�X7��9��!�w��+�i����xi�7 -���6�1|>� Y���!F��݂��p�T���f!�*�2�j!��2 ��k�R���������ȧym�o^9���ۇ1��
��5��v��#9�o.�wE�i�-1t�eM�����DC��� �IMKS���Ǒ�/5�ب��"�q����M����:�F޺���E��F�f�v�*d�a:yZ �,���';;�>�2Qg2e�T}U�[BB���Y7$���צ���޴��u�� ҙ���ѵ��a�d#�MY��n�&V4]�z�j{�+,��pOr�R]d�9�3�
��WnX��؇�"�)�>�6�je���Z`1�@�*H�5��w������m��E"���u�,bj8�����`�P�p��Y��VQ��?7z��hs���p>�Ǧ~���y�E�vW����B�&lXY|���}���c�5�{P��OO� Cvrz5�������/#s5n��Z��Y�����F����-��0�]p�8���������
�U�.5��A�Y� �9�����w?O��(��`�����%��l��r�l��s�8�R�-��<��PT���fc�6�^>��[/��چk�҃�v�`q�|���o/�����k֥�U���O,sBg�+�B�1f8��v^ze�<>�z�����H�8�O���K��q��X��gQL}k��	����9�O<K�x�u�K �:�[�I*�y8��0֨=DX4���K��{���?iK#�Si4��I�@)�]mU��q-���]����$Jp��׃�s�4�'�����RI�ᯑ��W�Sj1��ۺ�xDX`�O4m�ˀ4{>x;]'�ZJ �>���������"��۝�7dɡ���F�!��`�pN�V��E͉�����H�[����%�#8���.��^픾3�-�
Y�7�A��`�Ѕ��Y3cGc�ϧ���u�4x���3�U3��� ��l�(v��5��: �v��J�����ׅ����4�Sm&F}z@�7�|���M���[뀜����p]���Y�W�E��T@j^D/�A#yvX�������]�F�&��*�->�@ޯ���Z�d�>%�C��A������%K���T�1y����eg �KW�2?���|[c=��YJp�B n�k�^�<_�bY�b�]Z����Rz~:0X�r����I0N1/|�5s��\�;�T��+ ���',�mw��_��T)�
{.Vd.���#����G�7��'��U4�2}F����nyH� �D��t�O�Ij��k���7�	��|tT�C/����G������QJ3�g��{��]@>�^� �$�O��	o;��<�0R�q��'L���gj�U��K�n�5��ܐ�ى�G�1h����3���S����j~���_\|�qm�
JQrXJ�m?�Y~휤uԍ��ֈ�w<�N����q��vɦ J�cjQ�o�ciң�w�~[y�]���}G����r�v��
�/r���n�t� ,)˓aʝ�2Ѿ�~��!�=��J��`M�O���xlQ�*@�����"+���K�^6��ٓ��i	.��m��մ�tMz[�߇�Pa��m&�e�}���}�"'_k�����T�L!����`����]� A�����%��Z�<>K�O9��.r�t�j1�+쎎6�,���|gԴalU�(�'ٌ�p��`�k;W6ӽ�C��q ����N�A2*��(�:[���t~��Nq��Q�ӧy��O������~^�[�v|�@��$n��N�Xd�vvW�d\9f/&�N��M/�Y+,��px�a�q���8'��-I��~#����`�7�����_S�=�,c��]T�W+���jޜj�o�a�B�k|6�k��]ڕ����Zބ�P�����:K�p�L(:�r��4,����C��:�2nZ��П���q�c�r�ƽӒ8~�ߔ��|���0�s��u���T&�'@�W�k��_l~�)3��p�O`�� �����ZA�� ��%Q~N���z�܏�b*���q� ?%�#H�ߟ�ؕV	߆�F;�%��!R[/t�i��T��^�;B��X<�Wm?	)�<I�@Ew0�w�>�1�o��0bs=�ޚ+�k���������a����!��8�ud��q[���v��Y����Z"�r��Y:�
��~��͏���2�@p���ߟN��:�'�W`)�Q�.y���{�=Y�p��o^�:�]1����ӂf"
R��6�6��.f��v��G[�0Q{�N'fr"R,-��s���IN�n��+{s]�	7�q����\Q��4�g4���Q��äX�����;f��搩��Nd��ك��Ҕ~��f�+'�	�����f:[O�)I^��=�>^�':ې7;�li��n��25d�X��h�^ɀc��7�yUe ��sU�>��������b��=�Z�D{W$4FT/n���t���ţ��c��v���|5���S��L_�x��5v�������|�%�HTr� 񌫎�s�,O�Y;��R4Ua��S�p4���_���øx&����N��45���b���Ig܂��� {���������4��#��w�,����Dz��r �9���C��ƽ��]:�g�Z5���6B���6���s��G�����X*�&� 3�;��W��Iv?�sط-��x����v��ה6J�I D�s���|W�~x`�	J���݌��i�-���V<Ałb�[�Z�ۿ�r;vk�@���(���҈�H��?��q5���/�e���SX�s,SQ���V�mI���H5�pE��;Ir�����yP0}�c,�64]��35x�H�F� )McS�*E�ʙ�	�C�+�j�+�˙!��f��0�?��>�#��s˘T��������,�ي�@h�W�V��y�U��M��g�iw�^��t�-T��oP`#u��46��g;��a�c:��Y�����#�-����;��k�����F�����3=cd�uŤ�N�nr��H��ߪY���΀�,ȅ)�X��D%Y%g�� N>�5�,�T���d�X�$FQ��%1�H��,l��SP>S���l��W�����VK�D�5�٦`��j�|��	������D��R�k��M�6)i���ρ�)bp�$�g<�"�k�S���=�ԅ��Y�&;z7���䤶$������",��1�1׃���%F����0�?�,���ˇ);h�|�e��Η�v�qU�Br8C��u5`8�1284s��w'R�5|�������X�U�hXL���0��T�R̊iQݏo�Jm�9
�"����v���|�n�"Hi�h���"��� ���m����3���%�V#�4��j�-���f<���-c O7`m���@^6��}�,Qx����36oq���,'mO#_�MZO)���;�.�Ef��t�8x�sj�#y=V�e�uFl��=�i���K4b�)&LG���S�=G�5R���zd����L��� XW�A�ً��ta�]<��;cNXSH;��3���p�O�Uf�ޘzu�-N���H�G:���H���'�<��J�L?�*�l@���|mtIWk�5}+���s3�]I�a��]B3�%�}��S�0���_R^���-1���
��O�|'&} �7�Q�g�37��oY�?y��2�7�L��A˹4І��^?�m�%TxDׂ���sFZO}K��W��ə��m� ���:Y	7��;F�岭��p{�lC���RN������@BV�eU��@*�W�r�D��
�zJ�?za�xD]�*�^������8��:�)����/�]�P��FnQX���G���`�|�oo�i\���U��� 	v�~kW��U|������](S}��y�%�=�R�s*Y�t]����Rl*�<��˘����k�k4@�Ԋ��9��	!H�]��>��Y舵��Ѕ�݁$M��� -�n�x���Ύ�c�ʺ��۬�������(?�� Z�,���UMj����A�.��'�8"��(���sК�V���f��y�X��Nc���mZ*�>}k�
�`m�iD��q�g�����S2f��tlj�X���v����T�'Ɇ�Pȟ6��Z�?�l}PS��^DTD��tA�tE��NDJ�K�E�
H	���"B�Az	������w����?����}w�}��}ߜ�2���~�n̗y�܄��O�������Nc��y�966�W
�k3#��.2��>]y��^�<r8 ��܆��(A�p���S�����;�g�4m��a%1���W����C��UX��+�rA���F7v��a�t��Ԋ y�oϮj�8�\s��΅4_a���/��d�vlVy��Z+����Ƈ�f7e�6N���U7�d���-U���R��cE-�!�q���B�z��ix�xP'�ဎp�}�&W;�8ɌD߶���dz=�ݮ[�4?V�F�RѬ�3�_�=�'Q���n1�I���^��8Z�D���m?9f+���<r���븮����U;��\�](�q����@T�����DH
Si���>W���.�S������|�y�5Y���9W���U��I��j����nO���6("L�z��������Y�㍘Q,�(`�-�#`64�+=��q
�m�zW"y�<DOW�uy�簡qǵ��W/vTVm6�{�R��J�u+=���J���[H���%�خ��?�~Mʋ�ݧar���B�Q]�zqwn�/t`����s��/�u�v��p�|J(�*z3U�*e�`b��(ҏ:�s�XW�^r'��l��֕p�l���i{��aj_>@�P��^F{�;$���ԔH�۞ސ�q�.�^���=����V�F���,Дc}/�c�=��դv�-y����]���׶_�ԗA| &J�w_�q��$4,<Rvd�Vep�:%*��t?\3���e�e��n���ݟ,�Xm�3�Y�>���3!0�:�(Aן�m���+�;4�S�a9��ܟ9k�U�7���,w�KJRe2�
�������͌�������Ɏ���Vm�W�M*�ҳ7�����ë7 뵴	Ѻ�p1�o����R17=��]�� �}�T����[�����/C�D���oc{h#'�,��y��⼖�q�V�4��["jR�����fG�����~c���{�l\�x��}Z��E<)˰�ofcV���7yKd�w@$��:F��)�SO��})��q�85�Th������v�r�N���5����GVW͝�L����`��1m�z��ѻ�����I=���������ɠg��7t����(��
\���� H�n-a�����1y��в��H>˥ؑ�)�+5�5P����`�}�]Z�	�[{q�+��z E{���xu�FAMt�i7�6�]�c����a��T�e�<��򣛣��y����qT�����Jfh@� x��<گE�D�M�6#Tt��E�����ͽ;��=rmr���O���|W�V��n��G��{:㇝��e�^�ʥKݾ�^�a{��W�drv��#�6ܿS�����1��u\��ӯ��P�e
t�$ ڞ�"hQN}Sq��ր�<^;�V�/g��ukP3���2��e���`R���8��U�]UX��W��qxM�`0�P���a`�T��T���z���Fs���JVQ��� �Q��G�f/�o��G��ɚ �)���'��_^k��V�f�cB"�a�B���;�0���t3� �p��yM���j�cv�R���>�s������t�׶�Ӕ�'��I�1O�n���3a)ޝj�����<�UK숎��ƭ�ژ��*_+�X4��$�S\5��n~�����]{��p�&�"K�K��NGm���+��I�M���"���F�j� eX���c�'�,�:5/��_V�U'U�߄��j�x �+r�2���P��0y:K�J���h�<��F��.��Z]q%�
\;;n��N/��Q+��鱠��}� ɬ9f�i���C���0���q��j��|NV�	�@�ߋ:�����χ�;P*�)H�f�l�S;TB-�\�׼�mTN-�����pB �������� ѭ��7����h��C��5�KI[AW��_Q�+��n���9j�5l������4���?��Ν������U�]��P��b7��ӟ���j�.�S�6˺��o�k�%�A�|�f@(|E%]�	�=M�~@�Dň����N���z�8�TU�k�b����w=�5ɺ:�P�1���!"��c�TD(��o3� /=^���l����ء���S��~��Tw�ӰU=�.!����5�LY����w����畩\�m�a���Mۼ�[
Ҟy��C�69�36�	A�oҭл���,�讐�N��w�k��J��9�������U?�zJ��Q��q7uw�A�
goWn���ׂ��p��ݦ��������(�Z;to�;a�ʩKV��B���l�҇��WQ������.u���W��1�����������CJݓ�n�uk8 �v&��~��^�	�����B��d�յ>����'���F�U|GQ�k)�9�0D��Ap�aJ*���0�d�+�L�p���9�L�Nr��@��#U�����J��Ϯ��O�Z�9��_ i� �ú���@��+�� ��w�&������Ε��oNV���tu��MN&����֐&Zg?ŏ�����n��z=sv�n[��w�l��U�?	�[�*���$��̑�Z�Tj��3"�X��O���	�5^����S!�O,O�R�]�!�rJ ��8�e�8�����O�}�w���$��=9_;�L��AE��uc�]����`��a�dI�H�;��Qz�W�j�Ӆ�d��
�X�r�}���CQ��Zr?}k�G�*����,?_�8!9�~u\���=�{��b�#¼p6LJ�n�~�t�Ȝ�UJ���JgU�H����e|���.>���T;�6�+���ά5�MQˮ�:����k��3j��B4����Ͻ�M^�~%�X��XJ�27�*�!�s�r|S��uՋl��[�y:\�{ZJV	ykq�2�1K����Ra?�hH91%Nư�g4U�ŷ�]u5�Q�~��>�����?[�a�ۦ^��k�dhs�p����ۢ�-��M
���7��C_A�Mℷ~�g-D)D[V^(b�'d��C?ܠ����˸:}�_�k��`K�;��X�+"�>������{����t�]��u�28YŪ�;��٤@��K�]�ߐi|�}v�g��{-NR�\b�,6�Z�$y2�EZ�8$Y�Z�و�N��4V�PL��*��WhBY�W���G�$��1z�G�8M!쩾��-�a5br�7�S�]Yg��A�+B'^�6�걗$:Yn�+�ӻ�$��pn� ��K�A3����繍���T��|\��fG,vB�g�HѭE1�	��N��1 :�}���c�����_o�Z�j��~� 7"o9�:�`���y���	|���_�n$�n3��}>8	�v�^�L�X�:�/��O��v�nmG��;�� V,l/�]��h�d�e���)�5!�>���J��g���9�D�������!�b�K�5��;���8�{�����c߇$�˵��.����0 �abq��s���b�m�����\�HЂrcv�V�n�H9D.�a�i���{<v�Uډ�56�E�މ�)c������uj�-B+��!��������&r�8��Y�&�~o�M>}�I�#JX<�%ɏ�?�F�ʍ�c:���������� v"C��T�M'�-�>a���v����*��&���!:�GM�ySܟ$w/q��p�6`u�0����$�ڼ�y|x��B"���E(�1rg���Kn���� lv%z��(b$�+�gz�������*��EI͋�g�	�zȼ��ެq�	�v��$��j���_�]*ڽ�ˈ]�*xU���Zs�!�y����:�x7I��oǠ��F�#`�R#�*��8dT{�B�9p�nLĦOҽC��f^P��C�D����Ta�n�w���wS��]zq�>g�qM?�nU�Lb��$]\�,�P+7p-r�*mc�V�qr�Jf�.���y�b�?Cud�����w�Z�s��;5�V���:���7�n��,j�c�w�e���[_�ؘ�"�*/��2��}��O�_��ue���tp�+O_pǿO1�A8B�$8��k���|�3n�B^Y��w{���J	)��o��.V��(HC'r��~�y�GS���Kߝy�&��7R����=�T �Q-�.uҩh�!�x�k������5.�Y�b �c����C��9�j^ɧG�~i��S��'y<M�9���"/>�"Z�zL�A��~=L�}!�WzHǁ�ς�~�� �OP5���<[����k���^�i����T-z�U )޹�����g�蔗��[�&��MOc)�mp����c�Ivi�cC�ڍT���'T<wܫ^�	SQ@S���P��`g�r�� �8H,���U��J�E�v�!#�������	۔T�P��+�*���(�_���kk��f��UB���hzW:�S�`M����V���@[�Ȳ��	@���x鈦����G"x=�l�q����%�8�"���c6�|��Z9-o���ڡ{OMZO��4	�L���	�Ƚ���ƵԶw`ѿb�w��
�@�W;K����%;�_��� �k�QNA���[R ^�J�哧zj�nA�~��������+\�a���WQk����xꌅ3)8}R�ILs���|ڡx����+�U��<9�#�lS	���Π��'�Q����x
����3~�x���Y9'�&U��A�>�N���VC�65�$�ֹ���%C��g}\�Ml��?8�TX'�f��|A�<��?O��G���;z����4C�SV>$�޴�Z��4�]���}�؛G����D	�BA�� R�a��ܓsA���NKWЄ���2mH�V���_g��um���Ĳ��Ϟ��1~o	�@�
|�N��F���P%��#l��q���	��X���ߊ�&Nk�����������)�SS`�"�'�Y^8�Ϟ���5y�������g4.�����o@����r����Q�f�\���'S�Y�YT��7�>���S�������'�`�o�I���NK��)U�s��;�y�`�@�����[��^����������Q��j�R���vI�]�<8�W��W�ݧ�_���=�,\c�1�q��:}�v���sCB�p�v�]H͡���ہWw��&9�{�i�k��¤f?�	oL��^u�»Q�n W�E2��u�����\�S����>�:����|-��]Xm�H�-�*�!줌AbS	/)?�������\�!�(}fI�(u�_.ڬv~��R)j�H��Y�d_�f�q�(<L��{�y���*V^@��,�'���e�2ﺠf�h�N���{3tk�pf�%� ����=�_�v|�S��˹	'��o7�?��/K���N�@{[Wm�}z�3��=�ҿ>���CH���M�N$�ΩY���W�J2(ϓف�MN�[o4�������iX�uqs&5_�B9��-5��'o��#���M���~]��ﰓ?������P�4 ���$���ө�Z��F�LI۠��E�PX������.��Zo��q�0��ζ,�e�^����Ճ3��>��Kq�?��/J]����;�nI��"Q���?����T�������W�@C8f�=*#������a��� !4��c�N8oE��I�x����9 Šwɰz��\!�U}���8ɄYy�����.){�yej�a�i�L�4�]�a�=�2��0���P�}y�v2FK�u���[,{9���̈́ەo� ��G�nƓ*U�ï����.SD�k�a����z�]�D�Y�X��87E7�g�R[�K�H�(u��r�]*��='JO�����mI�m+5�W4c-��h�F�9e��d^Aѣ�2�x�5��܌�e�/V!�0w�Ot�>����G�t�=�4|�N�֤b�� �����{�x�<1�=��Y_1:������u�G�f�`3Ъ!2H���I�&�� 1��֐�ת��h�z�R-�6���|p]��HV&��{��W����.���L���v�A����V��5g������bZ�M|oh��A}&Ng`T
J��Z���&���[��Pi�>�px?ql�@*b�]5�;y�M�T�-����~}�8Ģ��ȡ�ϝ������h���vL~���8$����
�]��IN��@ߍ��

I@���^]����MDef�';m/N4a��WB��QE�ZW�� f�����QT1B��Ewx��:㥛xk~�B=�eݷm�D�RP��E<:J�د��Q�ӽy�yw�Bp	�������vX렽;a�k��g/f꽲�|	��C�g\"�$�_ت��>Ceg��P��ɠ
w��;$�����>n� 9v����v�"q�EM���Z1�J�6������{�K�
,*!;a��:���2Ŋ]��tۡVb�,�
:�K��+4�52v�аqO��ۘC�Q{�ۼ�x�ٞn3�"��䬨h逥oo��g�3�W9��lhvL�}�3ҵƏ��I$;O#]�IF}u��ޥv%�p��(�u�ߑ>}��,҄���s�*���U�M⵹��{_��h�Sз�׺u�IV�E�Ďz�}'�<�,n��^7��Q-�&�`�qߪ���KKȟm�x�[,�"��`�����9���
[��n��嵁g�.�|���]�ߐgށ�N�����L��zj�����P����ӧ���E��L&!C�"G�XS�����&t�=����)|e	����w��
�{�_��r��+/�����\��nS�,k�O�4�u��]<�E4�cE%�a�%��P�66�C��Sh��[:��Dv!V��*c���1}I\������D٫ �c�����=@�������px|�d���sʞ�@c���u�s��&�~�4�.r�I��˱�%;uf����ϽǤ�2?D}�'�=�Ƶ���q"e"�~�����d�Y=��T�y�h�
�(�i?��[bq���>������3X(�vN�AV*���t�߇�x��(�u��_�ɣ��.�0=�W��Gbo*���\M�zK�����T�u�ׯ�d�u���ZW�.��Ѷ�SX��g��Yf+��t��r��f���u���{b$����A��m��&�A����s�tr85?����74�g͊�ji��#��Ch�V4�8��	�E�z��η�uT�4�m�g��rY�����4���~���`��A�;;��
�f��TuH"�#���F�@g��=��p�$e~��)!�����+il*6ʀ{����ʯl��i*�<5'$}_�?�&���F<�΢�]��h ��~�ʔG��%Y��#��I��+�R�ޚ�y��y��g�&�L�g�_O��I������'�֔1R��L���~��N�Μ{_:B4��-[����"'��U��.����6fx٢����܍&��5���rBw���ۮd�5��L�6�{wU{��ֵ�iP^~��9��{��V�G����u�ʿ�-��2<\��k]�Ї���Els|N��g=:Uڪ��k�b�r)�D�TP���5Ie�1���b[�<|3(\���.R�$�	<f����䒛7.��\}�;S:���fzgס�BZK�jd�w1�09��i7b�0���'����EN�g#D�ɋ�WQ�Q,s��*�+�����@��<�ȫ�;3}���|�h��
�[��$�x-pn<ԡ�Br�5�&8?%��>��5E���mb�|3�"�T�/_׶�|��~]��yҩr�UYB��_M�f b̰u�hQ��=�J�G�hر���ڻ�	�Ľ�:C��������J���3࿟�><�	p�:�NN>��T�dq[�!:a{W�I2u%�Z��{��8�c��VC����j����W�b�����Y�o������Ѐ�K�fU5Fʠ�&��~��G�-ƘD�f�+���\V1�-S�Y����GZ��Tc�L�Z񘯌Ij�W����r��컴��x��|jJrD7�H�P"���0d{�t��	���뿮��<6>:#�!hcg:�lӴ"!�l���`�׍/N�$�� A���w��J~d%1�<����-1V܅`�B�>�ȫ��2�7)���-����S���3m�ZlDu��fώ)����+]�_�筽�粁���⭛��K�TSy܇5�g��`�[��Un��� ��nV�ϪD6�tf���c�@�k�- b�^���{��հlY?�A��,�epw�s���WQ���}�=;5B�헛n���5<_�b�2V{�M�`ab�Ķ5̔ͼ�(��ҒY�b��6�W���t�	�!8��a��]�d��Y?$X�Ě��o~�a�eiu�����M�� ��QQ��W�o�z���t�:�^��H���s�j��ڰ�r��‪¬���ɃgyKNQZK�f��t���3�����훠f�r-�8�߼_<^�޶���֭ͪ �X��)�����ՙ���4�+�	K�����Cfݢl=瞦���:�	��=\X�E;���]c]���c�Q�|��Wηnj��7�)j�I
s)�xZ�c*.�Ӹ+g�
��&g��I��]�������
��QO������ʃ�O�:b��� ��b?fMN���9���QW;�����\KJ��Jc��L�~"�JY����ʗ�U,�k7�kϒ���xLc�B\�}�`Ӷ�a��:ɾ;���G
^�M���yl)<��Ĕ��;�ڀOŦL.9�t�M�m�/���]��.�,�0�V�^�GR|��C5V�D�
�-���P"8�S
r��{��\�D����w�/��\�2"e�v	(��h��YÂ���@��n��xB�Y"Ni� LuO߳a�-��Ѓ���ΊQf�*o7P��=��E, ���;,T25��H1�������o�І۵
r/�_��?����-Pj�ŏ�zݛ�zN��韜�˻��+&qה�C+��0\IF�T����@�0?Y�E�w�������x���]��)9~��kD%�=������㥛/�"�a�.Ԥ�REE�E�	3��tQ�|@4�@ൕj�/.���l$����b7�CV��U�}�&n}ٻ�Y�?�Də���N栾y�E�v 6鼤�3��t+]��[]c� ���-���݈�I����2:[HGK�_����f�1��:�r<�1�jӭ��2�� �g*�3/>��}Ě���"����P��M���<�@��?^6J���Qr6J��6��h�mP�؝�0vE�ɚ"�������F>XUR�jh�����%�Ϥ��]��n��,R�43�����@%C�Dz]!$ R���H�g�����TJ�ՃMd�כm[9{��*�5d�@ng�}��Ȓ�ƙ��wfX4��o��<�h;����/U^'���o>�GC	��b��ސ퐢�e�m�BO��,�\YTa�ߧ��� ���s`�����1��t��Կ�h�}eY�Q�} J��f����a��+�n,SVz�����	�A����ns)���5��X�x)A��4	���ɲ�Sқ����:���T�q�q�����X�l�'�cL�Q��~�cުɐub:�:�YD���@�	�M>����y{}�L��h��!��Z��Ħ&e�7�����u���{�П� �V�zO{Y?2GD�^�j��P���/��L�Lл1���(�Kv��+=�)su'�in抆O��&�e����
h�Ŗ_����/9[�y8L��.�Cv��Z��6�R�ݑ��fr��%F],In��Rg�<���C�l
�рK^��=�Wc}H�r`�A[+5���ҿ�猴&ƺ=�Iq�]����<9�Ѫ�b���J�-�I560�a�LP������mC���l�y�[��tJ� �Tb�	r��ܳt�
��@��y@�C��	2[�.�W5��.��uW�L�E�ǐ���1w=f��5ݧp��<�v����<�e�YeY��]7��p�G�~O�<��aiLQ�&.wx��Y�Bx 1���a���ߠ�����$��w).�E���n��5�'��Ѥ��Ay���m{�U5\R�Y���������� P����26R'B��g1�5ٚ�3h#2T��j�Y�.��>>QI6+�
%��E��P����T�\
L��i�2�p	9�������O���*�F%4�	�:�)��w�vo�~�Z�V|�{K�Z2J���K�߄��h\��Eb��_�+�S��Z��%�G�k�aa�iiMCOO�5��Mk�F�Sҿ˕taK��i�;�q�����$��dq[(����/fL���Ո�p]iϒ�ՠ��]��R
��#��OA=G��N!���%��>I�y����{�H�Qu�f�6��H���	[�a9�8&=8�?O*D���d���C��J@�rHSy����Z�X��Ե9��|9�%"�d�ޯ�!�L�'�qg���V���Rԥs�a)xyd��U�O��b���~Ȍ��4"I>| 4�dof՚��e����wl�Cß�d�K�_��M��^:9��t3μ��"���f�˭�>���MF�ɒL�w�$�9wt_�f��(�m x���J@r����>h�"��V���E-5�����B��Me�����4< ���F�%J�+�+��o��M�˗I��5f1R�/ ���c�:��@	h����r�K����
��Z����`=�YkT��pޱ9 A�!�@�:��_�x�4��f��؁P ��VRB��T�ҿ.�#y�ɔu�?&�J7ui�'Kϼ�T�z�P�O��ڮ�@|�Q`�Z9k�@�᧝Ǚ2x�6Wvͭ����
,˖mf� �a.�r���{�M�f�&1�����;w%Ō\�х�2�w�XI�Y�Ѡ�g#Wz@��ҍ�w��c�7�@d�.�����Ql�C�z�s�pH�k���2W�'���R��\��h�/��<?H�S���Y:[DU�Ī?-����|�?}愦,j偅�Lƚ<��C�-
dQw�-z�Ai��Z[ĘǨ#��څ>����u���M���*�@���[��֏r�~�~������F4�_�QBgR�e�a���_b��Wa��A��U���]�׎6Z��-D�C�4��B�؁��~�����t�s�BKZ@X��ݪ	a}�(ҫ��,��G��3��NOᏣXF���F2��Z����}�b��I�\��C���I�'���A��+&����K��2�����u w�k77��yC��!sjvO�1�H#0E�q�k��s�隴����kr�4e�+�5#9�骬L|t���F�g�%���	�Ǥ��uv�v���8��I7�r�8��w[\�K�:�,w}����X��5�/;���H���q5���{BC{�"����{��T��g��,�q�J�fl��r(������j^�3��_�自��y+f9�.����,З,�[�u:1K~7zA�sw��-�tyqDCٮ��,����7~��XC��߮���]��+��X��R��ڜ�H��{ct��}X�c�ʍ�k����;��'3	��ip� ē�Ղՙ��w����}��b�*������
#"����Lʰ;�*Y:�f�, WiU"�%�e!��ym')�g���h�p�~�.�iq���?����#󘶥z�e�Wԡ��@KL��\��%Ft|��f5l0#��f"PZ�6iz�u�bXA����f�P� "^��	B<��=�e�1#d����1�+�e@e�gi_Ŝ�7K����K��r���H�u�M�����Ӝ����0�;"d4+�����|6��p���j\���s�o�ݗF��u�)�l&G���e7���G�N|,ss��x[��2@�%��±Bv7���ᓤ��B��"�''wÌ�N"mg�]Z$�`}���K�R�.�;jY���FmK�x��Y_��R�� isBs3o��=1�%���:~�Q)g\����_so�O@�F���6�gLp�-f�l7ǧ����^����m"�hW���H�_��D���zx���QhW��8������1��0 P\�qA��#r�^����N�Q~fhe7�.M�y�z����0Gu����A������7��D�y4��R�=S�O�wh�2�~���W"�S$�G�AҜg
�-�:�y�[I���޻V}�'S�Ҙ-s�^��VX`��!�2��������YW1y*�k��k*|h�5�?&J(��tp��)�U�ߡ/�|�d�42��V�9���?>��]��*t0�S@]'f��4�>	�	A�G[�Y�$��sp�<t}�7�'�-6eq[�,�0z�Q5֠�.�;g_����J����4-oI�h��!�G�}���a����`N�X�������gPb�m8#�L��̧��?R�f����p��U�z�i��FO]0��BΙ�тТ�2����7I/�5��%}A�y��`G�����]w����Ɓ?��\�_��Tʾ��v�u����n��B7�	6�2P�-=xq����u���z��0�G�<�������~ѐ,s2��^�Ru��=����nK�k����N��gn���*ع����@�b�.���������DJ���K��vwK=W�(��i������Mo-�(��:��|�#�t�~u'�Sj���e��|��kCd���I&�l�ݢ^��<��z�X!���n ����Ud'�q,��ʩ�K����;Ȱ����5q�M�<2�5#���q������@�)ya~g������/}�� ��o����f5��[z�
�'���ϼ���f�[?���������o�c����K?�XX��j��4���y^}�(���;�@!���R��ތͥk��H�|�q[�|V����PYG�j�P��{/}�:�dJܾ��,pu��2����)&Θ$쩅��5r�V���j��ߠ�O�X�pB��7���%`W�p�����OC���5��gU�k�.�Sl��J���i�6��eY#�d�קI��������Ė�F���i�����,�����jr�I��i��M_KxF��{�^LįeoQ��*ݹ�l��,����
�����(�K�A���h<h���|�sj2�T����J-�Ƚ2�	������K��]���� *�:��߸ֳ1/� cU�����:���G��������Ew��Y3Z�����,��2����VVC'�t����IKĴ/ꍋˢR�C�u��2�71�l�׃ĪR�qf����G���͙�O���=(�ͼ�>@���w-��"�c�u�4x��t$��0S���uod�Bk��C��#�oAr׽A�*����3n70�e�˂�5�&)��fXc?� ~u�iܙ�SZV���oz�N����q�߂���h����W;ӑ����,�+�i5�K�"F>��x��n��R2��_(6?��E$�t�$�?s;�P��-Q"��
��*�Z�#����h�@^1��9ܧP�f61��&�~��o�}�·y�h<���)�J ��|�
��<��=Id���T�� �k�C�<yq����V_R`'=Vz#Ѡ�Jby���k��ýy��J7���CO�%\26^║I&N��;���v�8B�?�jY�9a~����F:���Bx:_����}�fĸd�ȟ&�c��wĵ\ț��s�k��`
T�e�ｓ���g7����͝
���u�N7q!�1���t��f���6�y�-z�2�N`Nk�, #����yJZ���d���W�2�&�@�:�hi���ᑭ��&3��7'K�����'�G�3aA?p@��q����i�:7�'�ȴ@��q�,6\ �m��-��:�E5����u�z�Ie�ڢTd(���;t���o}O���g��s�<��[�����ok�Ɍ��M�ʳ� 4GA4���E�Uە��ߟL�R(�됭���fL������z��N|T�{0b.�'����C����ү�q�E�}�cS���6�I�<��6��.�"*��r�x�\��/HL������0���������e�Dޅ@�&bl?Q �D�������@��O�L�g�Y��K�z}�+�.c2K�4��F1y��/�+!����o�D
�X�!�P��z�bJiO�!�&��&g����T������̟�&��-�q�h�	ݠ����j�ĉGK���ף�A�t�ϔ�^����;=�]
/w@��}���Օ��޵����P7��5�8�˅$g�N�h�p�G�.D��	������D�P�>��i��b�긭��L�2��;�J�b����P����?F7ìS=�٣�W�Tp�I�z��ړ��4zv�-���21(��~�Y�p`���4{
�V �V�<�����aV�?�y6�P�*�"$|�sE�m�2��0�78�7ų���_��#`��Jή�,�-(����=3Y�䥲Y��j��O�M�R(��"���/�c�坺8eE@L��Uڿ:�'CU�x��չJ��y<�Ǹ~f�8�ul�Lvx��E@�����'��O�l�_�����8�;�=8A$4|n<���"�@�;��|��3/R@��Bw��3Ě����L�6x �$�]�����X��}g������»�8���㙩鷯��+N5�:�Np��	�;t%�-�/?H7��i�W��Z��H�����c�c��#�)�Ⱥ���a�+�E�����p��@���Z�����(���t�N�n>��Y��S7�4u�`�TV�7��� ���_$�՟��fL�*|�"��ֿ�Җ�Z�T�������?Ś�f����i��(��PU5'A:#����'t�7����;�L髱�M�2�uJU��ܝq8� ���U�͚��q�E^��Jէ� �/�����C�,�2�;�0��X��Z�,&Y�6�� ������4����9`ҹ&���=���v��'���|	������f�]�xg�6d}&������]�s���l6�ڪ�G=�|C�¹����ڬh��f7Jh�PO�9�ػ��L�KXR5����G/<�>�94����{+�.V�8��V����߯���{q=����Zueoo�$�v�h]����b���	E��]MЎ0��3~��\���������7��<��}�����FG��2��F�j{����T�}�fJ��c��籲���rSօ�4�F[�]� ��:^X�Ӓ7և֎���ʵ�w���b��r%�^Vk�[t�O��F�{|��'��6j���u���y矿Rg�	�I�3��`��~���5u(P���.���;������?�?x>����:mc=R�Q�e@��mpġ
e����f�'�hRn�<[%�FQx`U�ɩV��R�뽗�&O�%�4�[g;��^���)d��3F����*�+���,9���v����	���G���Y]0g�j���8�d~����F����������Ҋh�>��}��f[g���<J��0u=���O�|g�F�������w��̺��q�G튄�e�|c[�Yx���e���� ��3r����L���#�Þ@��ЅZ�?�U熫��Pi7Y���i�i
� O8QMF/��[����=�w4rX��~�A�J	}6h�gk񣡍����#]G���������G��I��� �y�W��]�u)��&)��;���Be�h�$QǠ���h2ߖL��*��/����L�p�Ef��(��Q�,�r�Y\�^�q�]]!R�w5��F��$�=�n�d�����&@��	m����#g��t�+�^�?5�#�[�3������=�6�s��L@��eq}0��RQ�5������@$I��S�����C�PB�.���E��ė2�q�������6���E}�NE���Y
!HO�n�$N{X��`z��^=X�tR֘f�Sҿ�b�|aB�L"�W.Cd��SQ���ӛ��
��՚6������1�DE5��9�@ZtrY#v�f7e�Y���xN�ݗ�¶�rW$��8�r������Ӻ���.�T��XuU�"��9�ww��S��P���~�T�� ��g�'��ӯ�M��C)�2�G�S�u��1]��TB*+h�4��X21�S���=�Fޗ�ٯ&����(���� �J�7^�>r�*�;ڹ�u��k�n8+���fg�p�ya��� ��]�����:2�
%�=גW̶��i�~��K���h��h���kM������^���e� ��)��/����[���T
Q}fa�zKeC����i���ɧۃG7Ÿ�
��W��?�곣�i~H��υ@��-!a����v�ĦN뽂�S�v� ���&�Mq�� mUV��?�UX��g����?�`����l̋��!�w���2�A�^��h�/�,��P��Y�#�]�k�7 �����7�{�l��শ�3 T�x%p�3	0���2�����gE�����nE�"���G�%�M%:o��:��D��v�Jvߺ^��m�X�o$��2��H�
\�\�2�-a�O�09��)�}�Lp�4��M+�iB��-dt�G=��z��+��0��7���5	�A�:���ve.�UҸ����a��}�N������o�m�:��7Φ���}���~��ȨQ,/��&=z��������s��V-V���O��'D��q�c����ɳ� q}�d��U��p2�+�_8���{��`�^s̺�dm{ܶ%ڡ4������WW�E	��g������M���6ㅨ�Bu��Ҕzn�{�q�U'�f|�F��J����ǘ)�+d~�=m��#�� Z"�T2�"�'�ׯ�`<5ItRj�R�G�}�'�s��O]cs_P�0���rq���~��EZ���J���'����-ښ����r!�V
�8~��)F!�J�6Ʃ�� ���M���zo��lx�U� ��x3ӵ{������U'������گfk�Z_�oՍ	��h�;#�c�K��f��Q�PM�����RI��F@�EJ�D�ADJ��K@I	�n-��%'Lr�Fm���������Y=�9�u���z��;v;�����ϕL+ߋM��f$�}������+�=��l9t*����w��F�ɼT�l6V7����^7�(U7��s�/���+6�ӷ���a%�нf*���ȯ�??�]����|��s=��u2����)�	�Z�"j�:ju�f�
�g
@��Mnt'2zg�6�x�M�KN�p?4��n�e��:�b9E���E��_����gk��hK��'�u_��%���T�War���IfB�}b'"p=B��sv��+������N�|欈����>=��|m��"��Z��a?��ud�ǐs]�������.��S`>��`�[ �o��zS �I�w�R84t��*����5�U��k�,�2�B�p���]\�ㆸ��a/��|�Af1[�*��d.�$�]C��5� ��Ŧ�@P���l|�qڣ{��]i��-�kd�r:��V��mLʄ��L��-�$����3�/�Aŋ���f��$��B_��W���1�"�Y1.d�VeS��,�2p��S�����{�Z�A�m?{��Ѹ�>40[m��s&�"3����M�ϒ=[Gy��3�����v�O�R��>WVp�dW�:���**�{tSV��XMm-yF����c��%�"�`��4�J�S$U*.��1�7)�(�*��Cn,P�ao2�	�1�ު�����T�N����Ą��0^b��������rT\�Z]o��b�v�ZqIT�,����?�:�,��h��o�Cyv�M�
]��jQ1m4�ƜH�x�'�	�]F݋���K�T�Fӓ9F�f�$����Tb�*|f�d(�Њ>�3���#�B�,T����dO���w�'X�\�p�������q"7R O8�0k',Jg��玃���]���T�7}Ҽu�rl�c&���:U0P��ܦ0�aR�D�ξ�n��C_M�A%Cw�����V$������_�#�}�T\
R9�1��^tD��m��m�����=��vC�~W3�<~��M68�~�p���4���]��zoZ�$��~��v�D��&>`Uu@�^ �R���'�J�'jv4=<���Vc�r>��/PB*4�-E��Z�Q�]��w�k#ʢ�Z��c>��H�ң�-W��*�0�=w�������s�4֎��F���y/M�5���P巓�V�ڶ��i��=���&o��jR�L̀����`!�_�֌�RM��QO��Ö�[V&;�653
�������驘3M*���ԍ���O,���G#�/��
�ØK�fየBz�/t��ն�x�&2��9��Re�h��+b�L�h��>&M A�#K����n��\I�y>��e�*��b"-v�!��'�`����I�5�o���v�ME�rQɕ*�õ9p�����]�|��!�_����|E��{���Q���i#�H]p����L� {�ʺ*m6��CXᗍ�u����H�!A霮���~��&]�.���da(�\�4.H�m�' �����-���٣�)m R_-��R�H�l�ܳ>!��:r�n�yē��8���jb:�o�����������(؜�w1x}��s�5w���O~Ձ;E�LӮ�A�	vӖe�#\���\b�g�����Z�B�BH==�z�Ms��޵��>���	��}�l���ʲ�'#+/dv�`�fgG?��~��\�F�.5��J�3|*1���t����	d:;)�+.�mMm�;�/K����=���{v��*3sT�CsQB-�w���q�g���2Iz�%z���j�f��Y1�u/�� ��$��.�_��86�X�{��.�fΕ3;�֦��	`[s�̋�Vx?�)t{����8�����Z��ڃ�h��~�:92���@���@�����շڪ�Wm��6�g�%2-o�iN�[emr8s�EZ��[��z�|'�0�]�jk�\AZ��6K_�]���Pl	6���R��R}[d-��<��2V}���ųF츠S*��]jw����[wO�8��7�A����&�f�x����OO�3�#t�&��~�S�^s;���Ҫz||t������Y����
�e*����6t[�J�����,$�Z�L����m}�bl�Ja�`+��e��c�+�Y#/i�Ϩ���Ȯ����,H���76I�����zZ�|/��ǋ�_z��uB���_�"�wH�~6�ӱ�����C��uD� ���w�篚�y�'`�/K�����UHr�l�%�]����ICC�]7�S|��`|������Z�5�������G�ϳ)5S^K���tQ�����%PO����'��V��ԭ<5M���c��Ϝ��ɫw���B�o6C\�%jqȚ��}r�BLYE��չ�PF�� �ƲM�r�~�u/����x�3��P��f3��������@[���B�,�"�=y�/��	(��7�i����� ��1v��d ������%y��9Tc�?�o��\ʀ���x��z-&���,:�t<U���t��g��� E,�	�V�!+Qѳ!��S�H��|� Y�ݏF�2���y����=O�u�������u�'g��Ik���B��'��'��4���O�Ȯ��&��"����ֺ%\�2(��G`���nQ'9w����O����C�N���.�Ϯl]�0���&Q��kwl�ޝ�VT�%�˺�!'Q
h=�T��f�#}4�t���G�u+7x���P6�
�&#eZL�=-��|t����r��!J�rm`%<�{�!�Z3yalA(-V�t��c�#*�|�Gx:����zi:e���a^���Rgw��)U|�8HX�"֞{������
 "h���������=��R�RV�����#�M#Z��ڧ���^XP-�U�(��dΊ!�p������=��^{�3��.��77oq� 
���[�m��c��8��:�#�L2~��\��:��%\��>-��1���Y��p�Iq���Dt�FYU�~W�!�c@�)h�2þ���R8(ڜo�i�Y���\��fǸ�w��d�=��`�<M%~j��(�|��9��YT�Q�<)9^�����:l�������>��ܸÿZK1�/�MD�n����-�<�FC5]��u�g��-pz��ѩ�@����F��{��-p0�����E���5&�n`<>�[r-�/��&���ı*f}/��%X����q�<4��EŶ����,����,	^-���� 4�k�*��ة)���1�~�a���5�M-9���r�(�������q�҂�ը�S��z?i���������JS�?��~��4�iӊ��s��<(ziB�n_��p4ޅ y�Ϥ<W�L�wm��O�I��bҾDXOM�Bі)�7ώ1�77N��BC�ը����;q��QU�u/���]cOW6�,a���߉W/�����K0d(��hb�(}pw��Ëc��
��x��O~���R��ݹNR~�pM��Qw�OA�_Ofb҅��^��0��1�%�!���K�����L;��8����D9�-@!{oꉻ���̤r�p�%��m�)��-�um��:���U�C��;�QsW�I^5�P�������x	�D�����Oo��y�[y��|M`7{ZX�aǝJ��'ys�逸�ycCO5%�
�'gk��U�F�[#�tx���i�5C��������z�#jcׂ'�u�G��B�޿Q�H&�����蝖Hp��s��w�Ns
<W�,��%���d��ޣ�GEw��ڮ���%EY�Z|��C�^���Z����@�J�_b�KtEE��It��7Wx]iZzu"=�-�v~����u�ZQ�����J��u@7;bر�e-H�m�����'w:�%�B�G`ka�Q�sH�Y�W���?a�A��^��٫t�/��"�c!�qT���o�����ы�*�*v��(�T·����ד�&M�+�چt?ר�+膒4��*����&95�
�;YvV���L���Ƅ
�1�|���{��\/I0����s��yވ�i
|O�v&.Е�*�ܛ4)�'w?�h��y��8}��x{�OS�y�N�K�O**���d]��w���&�>�]-�Ж��a�B!��uk]'�\8=gC�<�5�yN	{/���&J��ʵ�
�U�΃� G�Y\�Ш�'�G�=�1�}lbn$�_�Y�0��H����w	�Ou�X�+�@�(�ԃP�ݭ	��e|Ry[��j)<�Y��g�敩ԵN��">0d����3�d��t >)�g�����R���>�^N��b���׬S�M��@����*>Td'86�s��j�t�%n���xN��k����}�:N���*���Q0��Z��
��Y��������#���ʢ7�?��6��I�M���0�?)��߬FߵPy�F*>��w��7�ğ�%��T�3ߍ��0����k�w�u� ��8Qkc��GX�uB2F�Q���W�(h���zx�{���C�;�4ծ	�H�o�eʞ�y���㷍y]{{�  �)���h�a���뗾�	[S�+!�6��(�@$���W�L&�i�b[�NlYkǇ ߍ�Z�K�����'?H�k{���0�:Y������6T{������N, ��M�4�^T�=ky��̌���}��[� S�;�h���]N�Hhm>���O��o�������ڬ�F�p��!�s�a�=�|�5u��Wt]@���}���� ��\��v��|��5��T��^
�9��qMu�
3˼��vt�uOmϊ��VV����9���e����d5߹
~�"N�e�s�P������S1��V�i�bO�k��>�������3\T��_�]T|�*v9�Uz*���b`�G'�{�}�<
��q�L���ڧ_e2	��WK�]S30����Se�٭5���VՠB�����A����+���4�"�U�.��P��3��T��0�a�NP@��U�7?W�K�On�>�ͮ�k1� ���1�Ą�h�4 i�m�W+�тR��T8�;,�D��
7�ޞ��0�(p�3�F�Mr�ך��'��|!V�(dVm1�ǫ1��g\�${gLP'<j���Z�Fg8��*�� �2]]N��lI��AMA��lL;?��*���a*��F�8o���[�~���JVV0�A�=�9Z}3�(0�'$J���Z�(���&vЭ��X0� k�5<OMxo����{�:�T�����^���/�*�A����j��s���eb�s�g���ُ0�������;i�]-:˳�w���>����G�~s����nW�"Y�Ī�w)K��[�j��QQ�5�H����Q� 2�谌�hzWb&�&��	�bQ4%R�s���v��*��f�ѩ����B�>;��<E ��YF��c��FN��ҧ�n��b��ʡ�st����h�HI�n'����$�3���pP@4L8��H���M����mO������2[��G<�oTw����;�ٝerU%\|:v�פ�j?>�,A2�M#�d#�6�؛K4��d Y,H\�&���\؋�FV�>�!'�ɏby���c�3=��lI�5_������#��.QB�<��0D�}t[�*�2e����;n�w�B��^u�=�����jF���|��K)W�d��.!���F�F��*J�l���x�ͫʲ�Gy��ɤ艆[��h�澦B{����M".I�󗼻�F �����'0>u-_���#����HE��UA�*},Y6�z��n��,�&���%{�*\���.�+�3�3j��M�ޙH��~皬�mf>9�6������/��9��K�3�\��@!�����FU�k���U|�u���2�|\�+���Lˀ�۠�fٸ�C��=
�\}f2G�{��P���X�rX�6�p1�L�+\I&WIf:*���Yu,��Q1�N{(�rE�)"#��e��~L�t���_�3���� ���}���e�gD���W�̽�Z)��#��o��݀(��ߡ&*�2�[h�1D8�w먀���?2MÊ�\��	��\��z�jI��؋X�Z]�XWU��ۂ��b6v�y������	B����w�4&�،��H�O�x��Q�,�z��_�����"���~�Uy��v�Bx�k�9�(�٧�.��9qP�+=�˧&�;<��|m9՘�]����K��ei)����GE��u���t���^�v9�Sƃ��+R�{��e��%,|BIk�4n��(�x�m8A�,-9�7:�&:.�@�L��09��F��[�U�>�9�wE{��I]�}okzll�H�R�)��]_waok
�AX#����R#����u�ɩ����o��n}�h�}�����~�D��:s����BK�s.���73��yF3��� :I� ��+���SJ�F�
�e-f��?�A�H�[J��������U����̋g�ʪCWK��D�f�:�d���"��h�G��/.3�]���y��8}�%+sko>�n;�u�Q��W@�&z�yU��1�zq��蜽�*���d���cJ�+�I�wi�#Ъ�^�i�_�ҵ+
�U?ƾNF�� i Ni�i���y�g�k�Ӵ�賜���-�M������d�����1,�0�[A�H��5����I���)�O �9ǲ�Yet��	4�������)rX�IJ*�f����U�o¯��;��C�h�P�Qm���|�p���L]D�>�D��K����躌L��k����&Z����<�xW�*�
r~��^X�7Q��c���g&c�H�c��]�D�x�~F�b5m��U�j�O�x�=����h�ucK�����pK���?iį�� wc_,x�[ܭ�F�����H^!�}k������M��� �]�a�4�jd�����GQ�*(m�{Cο�V��;;[±句��e�������f��黡j�/{? /��6 ��L��P(��1�Yڣc�@��U�¿jܭE������˖k���aY\^dO�R���5�x��n�4I��Sft�`5:��N�ت�&O�O���F�6^p�˴袆�����v?����G��+_BB�;;�_�)Z�8�,�����ؖ��-���4<��[����v����У�k�%����@�[6-�a��:H��c�ʻd0���o.e���0�������� �c��	PF���m����2�Wp,��h�1�`l��e�}t��O��,�G���1܆�/�~4��w���^2	w�[�G/v�����N��q��Y�y�;����uY��f�&�Y���q�w�w:V+[�}7KI���D��U9Se�Ԉ���<�l���;�>׺N+ P=K/{$��_�>�`�ƻ�Fk��:Z�&��X�@��(Z��62�mk�-dp%��#����7�p��8��?�ub�:��f��a�dW�>b+�C��o &ź��.#7 �ۂBU�
��c��`���޷��v�lɧ2�1F0Oߟ��i�W�ޠZ����1�|��F�m�~�|�����b����*��0��kIum�n�����]�:�$yeXqe;U��X���9|��V���.�}6����i~�ż�d�z�=�����*{s�0�(*�l�f�hsU\7$%�Tqz��Z�݉��H��C�4�������Q�{gv�]v.k��hu9U,�zq��YF@p�wqE
���@�e��N�3+ڜ�o8Ֆrgg87�����cMP�Q1@C�,��砷
_��JK�r;��,mB�7�T
���9�Zx]czTF��8j$=*'$��}�nU<� ��?'��TT���a���N��f@ӯ�`�G����zي[�|��ixԪ�$h��/Ο���m/�_hVy��x�O�#on�����@L��s�rk�[��q��Co+�a��%L�p-Mn*��l�T��F?2��z�������*�!I��|��SΑ;��Ԃ�Ȥ%��_d���J��[ܾsl��yު7j���������c�SX�T�_�K��m5>�k�SWdk1DGrӼwrp�+)��tI���l����O ��ϲ+~ �0�,�����$B~��]�p9� �+2�t	~᪨�dG�g�=�I��
���~x蚮/��LR�δ^i����I��k�]�Q9#m��坝RPWX@t��r���'��G��P8���c�Np��Ih��C}>SE~��.h�=i#������X��Ee�qK���<ꓙ���	
��559��l�k�w賲�0F}j��Y���3��8��q|]Cd�.z���.ZBr��sh�h��>�|E��wc���c���Ӻ���đ�?���i�V3������Oe���.��]h�]��}�W��Ö�x�Fe)���<Q��C�%ĳ|�d�jg&o^'�������~�-ջt,�R��`�V')]�tI+�Y�XU�!���,����L �����>&Ԑs�MD�;�F��ta����I�2��R�H�V��71/�D�l������=m�vy�
�t�vm�t�[�\���8�|�&������k>�i��F9cS3AA.>�C�N��k�)��O�N��Q��˃�7[� ���⼸r��jy��;7@�n���ۮ��&�V	�U*���lI�²�\΢��j{�k�d�Y�G�l���E����-"dn�eԱ�9��`E w��L�5��B�ٳ۝"����e�@۝�GI�ְ�4�*�;���n��0�0O	�%z�>��&�����B�۪��買��q��U����N�10 ���~t�K"�*dBK�;N���
��PN\h-͆lf�q�\����_ˠ�:ʜ�M$Ĉ���'���W��0I��q�T�&<P�&'5��Ej��$2��ͮ��]�t��)R��Y����-?�tUH|�E�@���x�=
�V��KV8F��ɽ��88�Mw�?/���o�Z���u�G�!k�{�C�ϸ%��Q�D�_^�L����BͿ�j6��d�I,J*�ӻ�R/K�UT_8^�=L�c�6�mli����XF����,*�%�i��$��Q8Ϛv�Y�|͔k�vy�~^u��'n�2ޚY�kUW���~���\`�RDK�U�$�v���_�揷�W�:!@�~�%*�V��eX���"^��0��Qw[�F5�	���,�7.��l�E�M�.�+쟞uY����@�Ϭ�΂��fS.c2��fRϩ�7C��3���&�u�����w���Fɷ��p�<�\��ŏ;l�C��f/�8��̠0�q��ty�9������_G�.��g�ݵ{�L��So���i��mE�Xr=�*�a_��ą�LN���|{�~���Ryh�����G ���,��g�����0�����ߍ��C��9OE�X�6����Ҫ��{�4.� O9�輸���ywPz��>��T���'��ڟ�z7\�!�Le���mƨ��H�e���u�:������/Pa%�u��Q��S�9�[��6�آD��s���m%UgZ�ܖ0���\���و\U���V�ΝJ������:�E/�-������N���앎q"�[]��2?bBG�J���L�t����"eo�����eeL��=	Z�w~ilIQT���y��E�rݪ	����W������pY8��r�����ۤ&T~�r3jѝK6+Z#u^�cз�Y���n��S�E�����p��*eq�K੯��TK���m
,[����l>��S#��� o1-
�
�^���+���{�M�˯jȴu�L��=�<Z��.t)�@���A��LeX�a~!�36�@�Ġ�0s]E<��QNK�
G�'��k ��* \�hU{+�?�a��fD���$Wl��ɩ��|�Y������d���J:(Xs���J�������fY�ۯ���*ig�$-B��g( ��E�+C�>���C���~)(����~���&.���  ��n�B��7Q��L鵫/�~����'ϊ��L�	<�`"�6E�'����g=��ey�.���
{� ��> ��|o8��Qc�/�ǯW�LtpNsb�Kx��EnA�X��	���aӅ��Օ���1��A��î�T�ޮ�EE:_�/�ªo����Y�|�ݛ�A�6a�<�y��o{��Zv+	H�S:��/�l��'��w/H������>f���G�ή�w��(�������$�VW ��6�JP��ou��-Pg�u�����������髶::�|����̼(��-d�Ɍ�"��(�0����`� ��F��XWcYD*(�d��ˬ=�s�K������tI�jή�����ƭz��"��纕�	�
�.3���X8@�����GEB�{+�K�*B�gu��Z�=���r6�땔gi����5n>�:��o�v�=v��?����L֥uh��������¯��C��m��s����G����������3����U�dGGF�-��96�)V�Ϡ��^���>���� ��K�l� P�+#�p���B��U��W�1�FK]��gJ���L�-��Lv�� ][�,v����۫Q��A?�y�_	��;�X4��Dk��Z��	�U��V���m�to�D/^��p=>͐�zpT���4������.@mu��@dY�}�T���P1�eif���q��'�s�z�ò�Ĳx[(?��KP��maæ��Z��߂����  pdw�2@~-���Ӏ�b3/�qR����c�����{�o��i����to����	j�Z�l´K"a�/���%��c�mg�XhvO,��$�<����q`|������UU��n���LV�$0.����s����jk���N�_Yz�`��F��D,G������R݋Ak��;��d>�g����s�Pl�Ztz�au�Ir�NU���+���3���+��5��KO�����?�԰�͟P�a7�90ժ�h*P>�/�H�7�2��.��>���I�z���h����Tyr�|�z7Kk�NyYPP���r]��o,�T�a�,\�2yC�q?�����s���n�%�� V��nr�"��r��$�
�d�*k��jȖe�D1s�P��.t�����B ݐӍ˒b*���$����0�0�Pq�(_�uF�6 P@�J���f�ƫ�7^��΋�$��l�Ͻ�o�K�~��`��bO�3;,�T��GS���)Jl���m.&K�)F�8Ja'=�a�1���L�Qڥƙ���:�:��ABJd��I\g�0pUǷ�D���/�� �p_�&�f�(�]�\�>�l�4e��j`��,b�	0�!\6�PZ�����|���|��yP�kf�S�#gߓ!v3c�g��gB�c3�uWx�����.#�7��3@Hq��u  h���v�z�w;�?�ΒM�_���0_�90���k����ȯ�!�� �I1B<�[�h�ii��	�ޜ�u;a��u4%P��1���]��RA�.�J��=:�̒��={7��D��ڍ"�������G�l�ښ�0���Y�%u�m����e��3; ��eD?6[���!�����\/��ǐWcݎ�:�Mج����x[T�-w�뺵5N��(�o w�i��U׎z`F�^Pu)������C�Q}���ϟ��g�/��������R�!](�xc'��l�4����9F��m��Ը�ce���zF�֙�N�ʂ?���fA�H�����i�3U�n�3H�Dl��ɖv�ZjW��Ed`���VuLN�Ć����m$e��J��e�B �(�ޣ>t?\��Ĥk�?�T� �B�F�'{XC���&l ��W��.��+�3��N��a���`��$%��O�&����+�a�;H��2��3ɅF� "" `rL�Q�G�\`$�^��M�� ���6/��.#�T,U$O1���7V-�1��,<�^�rci�����Zb�<��@�����)�P[r�fo|A�u1!��O��2�.��Q���z�$�q��Rn� ��0��y�>��M�A3�m��
^�/B/�
��מ�Il1H2�Q����WU_MuZ������� �Lz(�mk@��}�S�Dt�v	5�^�Ӧ���g�oݻ<xqU�P$z���c/g��Ő&f����������j� @�[M�Rꐎ��X7�V����z����c�AVҪͰ�x�� Y��m[�JC���]1C�R��c�g$β> v������ϡ� �[�OKYېGo}�]��҉z<��Ж�=i�t�����0���ݰ�+���P�B���a)&���S�j�<*�)
�2�~�d�� k ���Jt���!��l��r����B��Qlg�!Ǔ���W��LM�[_��G���m�r�l���Z3�W  O��}�'�F������f+���ο*�l�����Xϭ�����im#���8P�g�K����,���Gzip��0�����ą�_��u܇l��B��_�T����&�]�֜U<+
��sh��Ϡ��;`A�_��J[�xV��lLh�,u}Wb
^�閳#l&�O9�ŷ˙N��iƲڔ]�Xy�x�mLر�o����Oː3]��na�����e�g�N��Y�G�AT��V�\�]և$��j}59>Ζ4��;�^�n~q���,\I��F!�2KS��ݟx�Dm�X怿}h7=	��
�����1�/^�!t�D�z�A����a�}�=7솋d�1'�+k1�������1���On<���0�Lt��`�^��|�q��<H�њ�!� �j�%e�� ��'^���b�Ѯ�rїJ�!~+��;�|�1�-8q4xNW��;�X�v�)���n1���ԦH�u��P���:����_�f�#dqڍI�L�p�W�A$ȜƦ�t�Gk������I�+��c��Т��6�u#���	Խ�5+�H��K�`j"H��W�%s���L�<������6*��I3�}K�ی�h.]z"�F���$`��:QJ相v�Y��� r���(�<��K��7�}]�$�������/�uVVFd���-N�XlWT�;c:^�K��!�r�[k��۟�M�6�L��(��FGU���4i����P@�Ķ��.,i�ۣ��e��3����^�����l���J�h�Nx���4?Y0D�\����%�G4���T���_�h6
0�ô��g����@��٭n�L֪_t���U5�0U��3"�6�*�,�����0�y`�w�/w����їAfG�Qcڍ6YnC����6 y1�Dz �HW�u�5�N��Z��J/�@�}�^t�'�٫�M�4� �j~�o*�v�Q'�A	��ZH�`KE�I	�Y���d
O�*�DE��mĄ�D�s��˾
I�8���Z_���yi�W>2w��7�D?�^�Xoo�2���}��[p'�,`.���۟�^��c]D%6�Ƌ�;���	o�\c-�Ͽtf	��sY��]<�~Y��J��,��<s��]�2�g/���ᕜ��\:fA�J[����iܿ����2�N���/[7-�47�gl������z}��|ɪ�z���o�K`���h��р��"�Z��4/Μ\�;����7pUXɄ
g#v�y��?�P��i���v�M��jѻc�"Dd�n�:��~�8�t�����v���8�yS���ߎ��J��V+���6�큗�q+����$�X !?O��(_��]�_�>%_�ޫ^:�A���I���Y����JM�R��w�
7Z�k	�F���v��n��{h��f�Ws#����T��F0ID]Q~Ƥڗ���a���5;$���FƬE��
�i�e�q;�-m�4o����W'��5�?���H��`�+oe�篧9<󞾹�*�3ǦF9�2K��މ���N�Y?��mD�*˽!z����:&N�f+�#%� ���yNL�$|P���dTS~Ǽ�: ���
RX����ҕ(���9ۃX!;WCdvk��V������]���'��.��;�kO�_�/IcI���L�<�/X��dt�%6򥬭�j[vo�=��a�&�R�Z����R3��x0r7P
9�W�猷���Kek^��i'>�	���$U���w��rF�h �\0��X6�d| �Z ����ha����=)@�"�JY��k/��? �9-mlU}e�f�����ɂ`�E�����e.�hF�zDB0�SGyH�32?����1\I��0���m@���׋���~� ����?�>$�������GmQ��=�
N�Q^������7���~�:�9gR���w��x�Mo��r���@��
r��a5�ٹ���o��X�n��q�K}�.3���γ��&)���M��nfYl�*��2�-�u-�Q;�(�Aj�P�2�?��W�Xe��Ac4�AF/QT;�BAɬ>�`Xsͤ�,mo�����l�� �x���ŗ�~�|�ܬ�J��DyT�=ZT��M`4�T��jv��[l���Bss�);&�,�I��zK��Z3���h��>��TqΔ1pG|��� �nmt7u�k��t��osG�T���5@��7���Mn�I�Y�!��ǝ��N�_z��(���T�M����0!�z�hy�C��
���"�Q˛y%u��:���Qƞ�"��S�h����o�}���E�mlz2�`�ٸ���:���l�*4�m�V:!��ٵ1*���odnF���Ղ�e�jҨm�ҚZ�����2�����V}s�n��l�(4���[���-��aB�i��V�%qg��;��~N[2L����}��<���QF�t�^E��L��6�a;���ɛ+�O��@KЖ�1�����~�H� y��&���'����"ǍSƬ�u��2���2C'�L��<:����mI��v�9���h�3MZ ����.Dj�^f�+Ե5���o�N�G�ofj�H�d��&�!�D������Fq�Xi�fX��,�r���8���+��-\ �ܴh���[�]{��G����plA w����C@�����>�e��c9���]�v[�1uB�B����cA'i���
J�
�It��r�a\r�:�:b� ���9�\X��ͬ������D����Xf2����QK�RA�책���� ���C��Ԩ�4��V��!q�U�[x-W0���ߙ�~B���nYc\�=��������a��{��ſr�1����RO�����#}�� �1\!���%���D\\9�*w�����������:��d��l[S����~�ڹ@��q����?��κ�Q�T�9�M�XOͰd�_�J�;���D����:Nن~�Gr�<����������7��g
�o�&�l���Z�`�h���j�!���;ů2t������"^� ����
��%+��%3`���蹯����}8�O�z��M?R���8���Y�{/�KZ���W�9W�5BA \��w��w�
�待;�gY��y?N(XB>\a-�W@n������v�1	M�HXV��&�?������a 51��<�6��`�l��f�$Y�*4���v$� Q"]�Ԍ�r����
�t䣞�{�����&��.�g8g�$W�4w�N/�p����ёE���<����23��~��9�2�S?�F/*�)�4���ot�A��f\�_y�`��8�ꭣ����l�gǨ�7�v���P�}x��c�t��+���y[ҰP;��U�?C��>��}��F��̆yh5�m��߽�
��iC��/7jK
�'_�T,��"��Yy����UN�����P��{�7�s±W�A%S���Hr3[�4�X:K��He�4ҪA�]ʙ*��$8�8F:$��u���ewш/~��|����3z֡h����%�%� S^S���R��������S���vZg)�_��E�DSX ���Lc�T�taV�Z�|C_����b��j�ÕC�=��Aj�]|�H���|Kk:�b�]n�(���X��а<�6?J���G�NEVM�On�^%A��b�굜�.˓ ��e	Axi�D���0�r`|#Zj;���p}�Q=FO���-�F�����YE��.�>-j�{�9y��9&\MYD��>p[��$oь*�yk������Ĭ�b�V ���xP�ة=�ך�	�]r3�oZ'#Q�M����cN���s�
x�C9�-o�.K��B�{�ڡ�b��1?I��N��!5]�鮭UTm��K��i�FS�<��J2���T�;m�q#���;���O��E������.���BGՉ���c�$�����4Q���Ԅ�@��Ոx�aZ��]Z���a#���N�Ͳ{	�{�)��QQ�5`Vޘ��6��ҡ��M�2���\�"3���E5�ut���r]X�n���(����_fU˝w�D~{=�mtL]��g
��D�d��$��&�ڭ!㺆S,￑�r=�=�]t�e�E���l�<�z�nJ1&z�˦��g=#>�>�9p�LU�m3$���m��ʴ�➭A���"$boȠs�����n$���������y���ݹ�V"@����̶����}�ױz���$VL��t��h��f���C���5���e�=�ߞ�[�r�Z%A1*�5��r�kgMcC��dm_�,�oe3�o���������{�p���oX
N5!� F�ED7z/ѻQ3jBD0��މ^� L�:D����:�39ϓs�/��ʇmf��^{��~��޹�o^��,�r���P�������=�9%��ؖ�ł�2v�J���g�`�{�oJy��Dj˼}9��t~ӳhXm֒���/���L�����ؔ<l\��I
ܒCL9Bxu�m��ſ�젛X�@��;	s���?Xs�$�id`��^��lWT�t��
ț�k�F*emS�y#Q�=[\�D+엷����|kH��M�W�ژjY��=bX9�	-3�vƌG
nw�唰��<��Xt<Ɯ�2����lt�mQ�5�C��>O���:�pǾa��^��u�6�r@�Y�iIG��F�0Ӧ�'�nE����:��R��/!�Y�Hv���2J�e���^!m�&��s�e�S�Gx�6]C�Xv+*�|)����i��~��{}�p����uļ���`3��I��cX);@�Sd�,��y���#2��e9ƁQ�%����Y[a���H�ZW�*����|��6'�
&%�b,h��I���G,م�=�~��	T���bNg�xV3J&�[bP��\?��ʓ�Ny��x�9nDg'xB��L3�� �-V b���C}a�c��*&;�G0DY0���P^���9��H1oN4m�z�X#�"�uځcl�53R�V�0�۩��[g�5�}N\����(�h��r+��}��'��K�h;�ԡ76��?���_Z#U,`q����=#�ӟN�*k�_����Uۇ7���<��٬��>��[50:� ��sm�䀘t�7"����V�����A�Z������P��{��"5rM0��H�y����^��$(C�5Ë5�:�g�����lFB��䒐��!@�����W)Jŏ�}�瓓��?�����yf:>3��M<�2N��$P��Tl�P�Q���)>)V����A.J`Mur/���1�:˶��|g��!.��꼜?5�������y-�U�=�{-�2�R�U��l���q63Z4���]���x%q������h	��m��r�˖�����R��,��`������ۓ�j�����Hno.�k����f-��̑{.U�e"�3kN���&��e ��W��V�a�1�g���5b- P��K+܄K�P2C4�������,S*��Ag[�Kp�6�IL��s�SMZ�K��q�3��f��&Z�����nr-���|�	�9�L��=�į���]省��m��I�ǲݡ��7�B�j�0��d���cng/��$�z���\U%H�.���_����&��*d�h����Β���hN{�f�\�컩[���u���ER���^�i�^�����UFy���,�)�Z�#d��/n���($�L>�|�UN���%���"�7����Bm0�A(&PmU�뾐�=���=�7��y�Y9��{�]�E��;�u\�� i�b��(_���"��<� |8���47^`qU����r�+�TX��v,8��EP�����3;%����f����i�A��ds^�3��t���u%#�.m(���q�f3��Q�>���GB��e]�u�q�z~�vq;�������IU?�*�p#����D�2��� �l���b�
�j/��w�����7P_瞰{���촩kX߄�{�-���< A��1��BK& &7a����M'��˗�z��$*J��.m9�؇DR�0��r�׾���-���)��ۜ��ɽ���~�j�@a9G������yv�E�f���Z����ȣ#;�:��Ģ��Ҡ�&�ӻk�subك��H�#�S���V�QBD�y�@���'���R�U��$�T��0�{��Q#�"�7�oIu������߂��k�/�*�̡k_c��S��]��D��a\Yq��1Ȏu;���er�͇��8�u���� ���a��Z	���M��/���tuD~�]��s�/^V���/�+=e���i� ?���}Α���`]����0"]#!�/t�.����/���_S������GI7K��=�)��P�'�K]�Lۻ���:�
�W���?S H�DȪ듃����_Y]��y���'�Ϛk���/�D{��~5�V�!7MT�����5�� �����ӌ׍���$c��e��>���m�����b�+�夽���en����!�~�I��P�'u�:-�����R3`n���A�j�d��S-��M_�����ny��%r�f�E���oԱ��o�r��;Ɓ�E4�$Ww=6ⅵ�9���gj=M-�R�B�6}�<��,�;�%Z&��z\�?41�ֱ�,%�s�E��`�|�Uj����9K*��%�.�� ���"�Ei�}�R���i]?u�ܛ�ԥ/j�=L!f��{V#���aO8ԧ��)���!��|��W�~�X�_Iru��~~W�KH2��	8�u�
��6�۱�jM��W~�0�X??�\�)�Y�r�Ɓ��l�T^}_=q.\���Bu�>�X�v���U�����v�ߎ�������tt<��c�}u��,�~�����Ӎ73"����ҩ�3;_E���Rb��j��C���>�G艳���B�(o?C�	s��aU~b���m�����������o�w}�;y<���uX�l5b��1��r��u�ϩ�
�@�L1
�	O�>v�i�S;�>7��ouo�qU�^B����!Ӕ��i�[��_/+��U[�Y[��5���A.�u����xL�}�_|��	�u?���E��Zu'k���K0���LK%�����Q��wNy��ٟ5�֋�<�O
v�8*8;��˜؈�
B�=}e$~a���fD f�|ۃ�]�8��E��|�,d��6�g���6�|���Q�ĉ;Y)>�f�*V���>|��PKQ��l:\Q��h�m�~ډ���4oG����ߟ�tֱl<~��Re��W���'�nؐ���Hs�f��қ�,8��H*)`��}�1�/���,��V�_}��V����3orKeL���E�G��	H�P>�_>M؍%���-Q7��^a��5X��qe���+� �2��nܝ �LD�\����粃����iP�[/�����f��(%�|d�pkIq���OcR�>DI���Jc)8nF��'EE��*e��J4ˁC3�L�s��5ę|-�l}�)�}��*��5bGf��$�P�LF��Uc����>�-��[��k�'��
����"3���ny�y�GI2�NQ;�>����S���NJO�������e��6x��[H�����<��6��x��g�i�|�M��!��}g2)���S�	�t� ����ٶ�>j�s�pp�y���������1EuuL�c�Ոx��Ϧ��D��y�'��b�x�_hb�[�I��HW)oe&�e^�4��E��������L��R'�^�Xy�e��њkVB���m�4�����7G�)���n=�|��=s&oR���ӊAU}��*s�ˏ����ó�;�>�C�+��<=��@p%���a����%��z;�Nʮx�@�,��J%~�wUJ��e�rX[����Cz3u�S���)dށw�DA�o<�.2��9;
�o�|+2�yk��kg:&�4�CO�s,%dEi�4Ŏm�o�}x35`�-@z�<Mq�}��*�7%}ߜ��I��ID�����R"���)���>_�%�]ޣ[��eA������U�l��,�3D����.���-���)Ju�R�N���d������w��C������32�O�B�������TL��}�b-��m�)�^ �#�e�R��'b�b݃nSH�}҄cXq��B2�kޤO�U]gyv}+��?J���T)v������Gw���˝�ߕ%b{X�;���:N�E}q�E�:B-����Ŷ�D~��S�ri�Ɖ�Q�2�����,Gui��3͈	��d�����=l��b:�L3H�������R%�%�Qޮ�� �sd���Ϣ�g2s1�P�k�Q��Y���e�]U_N��煈v]�)�[���E�4�E _Ԫ�\rC�4�D���0��E����얳g���FS�b�p2s�	�8��T��2��Y~j��WT�<��+�Ի��0x}�{��ӈ[�z��l0��ϩk�c����2�E��7�A��IUV7q�L��U�y��)D��u�m�����p�@Q�z�pm����먬��5�x?��L�s�di�"�)���2� ��0���s	/����9���q�M�N,�������jq���ݒ~ݤ�8�@*L�I'���S��t�{I�YM2eofe���5O��u�E���g���U#Mh� >S�\x��*d�]ZZ*���pSI̵᭠�?Ne�Ӟ%�d������c��%��
!ܜU�����*~D�[�s �ɝ2�k*���]�� ,�CFm�'�~��u�[MD0��Ƀ[��������Dȼx�j��
�B�0 d^U�|�)]V��bw�A�l�O2*1�I�^X�`_����%ހǢ�f���杸)�,��d[H$��;>�o��K:})c�#E{s�q7�<nTW�u�FVʚ'���_73$5�S�D���6�Vnu��Z�AZ�q�DM��#����̽��S�B���Ȯ�*��9֮2����x�D�
8!<F�sn�e���q�ݜն�qNK��l��+���p���lTUV��C��W0s�i�k�ĭ|�p`�d���X�?8HjA� �8�L�r~c�~7q����kb�;���߂�`�������hқ�Kl����f�l�2}��z����q�����-P�i��D2���x��(�T�XԨ�(�$���/d�jԘO�>?}��'�P����C�W���GbՃ��LϬYգ#)ހ}z�ŭ"﷋���S�azt�bV7���WQ4t����7Ԍ�*�!L'W	�3���q����bIT2W�R0��d���~���/�į��jvY��O������Y&�����z��/�lgs>BK��U'nR��཮.��_�>3N�+�o��<O�A�Y���tX�"V�o��m�ٍ�@��<b�*��PJ/�3_q��̋X�};��`"k����Y���Z�g����㵥�T�_���9�����Mҥ��4�A���Cɸs�ri�UFV�?����+8r$'U
�7�m����GF�Z�\��~��HhQ��3��_�RT�;e�+{fU�%�ӉAw�S���v�sGd�TV�G��[�M"	r_/�ݑ�<<=꟔v�n�i5ҧc���M;L����8]��Y�sbf64L�mh��x���@m�h�/`o��<�0��Q�i�����+��sSu`�l1�U��I����0�O���a�!���||a�`���TP�,R�j�jϸD#kH��e��K]D�g��'�w:tQ�˜\Y��̫%tFɰ�e&���J��<����	�ei	� �]e��!�!��xL�HpM���P' �Ⱦe�N�}�0��8ei0�.lbˑ�M�G(F�sy�P~��=-��M
�<�8����(���/#��:dfl��i+|a� ����ʋ��pxz<���ҕ2�J��^6�����s���0@%5���؀Oeɍї3�0��b������8��Z�0��� C���7u�M������|9�c)���ga��R�Ż��1�v��O �z�-�{�W''����˞B�:0x�&�Q��Bӆ��!�2�&�t{�7"�M��j�C�W���_���S��Rڂ��qkѾ���p`�cnH*�.�R�!���]"���v��8Dw�wn��Z�(��Щ�'��:�-	�3�Jm~�:����4�l:��e��X�]�1u��tD}��?E��I�X )`5�D��u��(�nX��ݰL�3՞�������D' �����JPr>����	���N�-#�԰}7vMy��I?�^F�#q��������#K�m��g;�B��&���G��	��סq"�Р��&�aMlQQ�	�_�j���e��]E��I�xq �d�L঻�Wn�-�����4EKFk��|�Nk��Jb�P\����0N�ю,@$m��ǡ=���-��f����M�Oq��\'�V�6xf��ᔋ��~jm�!��Αv��*A�T \��k$�tj����O��ƔŢ��L3�{o��!�Y�n�PPΌOW�U�>��:f�!E��a��2�(z95�<ŽV��@����{s�	�8b�2���;+��:�׶�0�ߴH�>�i����w.*;�!$gSd=�ә�ڍ{ʵKlm+�G��FI]���c�
��~����$]P�{�Ub)�ڈ��g�z��Β���*�95����qT�n0S���Ǯ�j]���UP26��?�Nl��	ʑ�/�oYʯJ[S�:Z*9:��?�J�*��NjK�/,��!���5H;��y?��lb^���hf�<<go�)�]�����5�]�k�0��-	�"7���V'Q
�/8"`>��R�7��
���Ą����B[��z�%�a�H��>�p�/
nH8����7!�-��&4�7L-�M�w[l���U$���(x�%Qj=V#!�Kp4��h{����h���`�ӕw/�X��4f:�@��u-�B�nEPՊMu��f�DV�7���9���uJ�{����,����'�IFG2�J׫����.��{EKvD���NF�]Q�ۯf������Ӛ|��*šAW��ݤ�ܤw�HS2�нj�dq�6_���E�ju	�s-8 ���0-98��3_�p�W,�up�2��;>݁:o�婒9MН�.�T�W��ދ�Xb�^���Mm�ud˄4��*�8��~��_�2�|`C�;�v�}^����n��*Ç�Q3<�=�:˥?��L@���>r�R��+���$[9-���r� l�1 �V�x��CeӅ%!� ^�!���9��o\Y+q���J:3��K��7]<.���3[�ZaL��$�V��|��B�MI H�!7���u�+׿�էF�h����+�d�ݪ��CGt'�}Z���KdV����X�E;u@Me�� `n��3HS��?�[�~ڬ��n�e��������_�)dD3A�
߮�s�C��\o�oTx�,(��ZʅoQ�8q�EIs[������>̫Q�����?^�K55�l'E�B�1�+�c�� A�mIX6�䬱���Xs-��Bl����� �d�jURXa��)y"��}.{nع�j�ڡdR���(l���x�VīH����%��4��T�p�^����=N.2�h+}��>h���&7�� CV���y���q~�����#Jk��t�C9�F�,���68�� p�\�����3^*�Z(/�L> ��╧�R�]%��m����n�L8oއ�K�U�13u�Îͯ]��ĽS�7���Fs�t�;��1U(=�Wi�W5Rg˷�n�8��熰f�8��Z�h�*��JN������6L���E_�7{�B�Hɨ;H�Sv�Tg��,x�&_�h(-zde�k�/W��PՖ�������\��2��`Qx�^5�� ��� �"����Tw�)ą�暓�\Z�,~��:��9xb�~#���ٌ磐�}����4��mɯ=��4�����TR{�c�ʱ��\�ڐ����������Q�O������jxVf�%`���i��X_�3��]j��������l�כ3(��]��"��! 9=vI3>�%���E�ӄ1����H+��$����B���H�Ś�M�0�z竾nɫ�3p��^}����ƺ�ҷ�vi�m}�NW��������U�i�L�=M�fw8�gd�,b�h`�A�=PR��z��xR�'�:���IB��r~���e��ݩ�$f��@[3��]$���I��L;�&r!�f�L��}51����V�̿��A������tU|gq���+�w�H�g�I��"���Y����tz��=̥��3��L~���r�qE�qQ2:IP��h)5�0_6���T@���<��˫��/�\Һ�96F�I��:�r��I�94�Vg'�c��!�����$D�ʙ��:_���0���Ȓv&�ElZ]o�5Nε��4��R�M6���T�Q:�9�%]��{x:�O%��o^-�aп�hB�DUn}�|3��Q�����ˇa#S������C�`��V�V�Ѕl{��~5�K�~�(��'��o�-A�Nj���������i�z�8��u�i�h������ҜV�~����r�T�����5���u�����&�ӯ���7�z6��g�������i�#�Ȣ�n���ܪ}RD�9�
y8v��K��\���p���nK+hJ��F;��G����^�T��"��ƌZ�B�Y��J�g �Ի�G���d7:)���ejw����N����ư�?*UY����j-vdg�+Ґ�-]e�6G������s�Tl�L�w5�Kg�a�,��94*�q�Dnמz)���ƲJ�@4a�ˎ.�͞�îFԌ��zd=wg/���/���t.)	���ޮ��/�󏒲U;S(�M=�Ҳ�:�9�̌����-�OT_;T~sb�����8(�,KL=���� Mm>n �g*�."`�J��o7�	B��Z[����z`��>�F��o���3�������v�q}����?��S�)h�����_��R���h=�5H�G�8��`�ZI����J�(�:iC�/�uz��ğJ���f� 1��V�Ieǁ�[$�Z�����̥%�)�"CY�-����Ϡ*��.�����Q~h�����WK(����'{�9w�&^D�l�`��_m>��I#��ՠ����v��M�+�q�ؖ�C��/P.m�ө�noУ7�-]~��	�R�M�q>��9w>k��O�B(jnN4�ZS%��G	F�Y<Ե�����^�f�1���&k���7pY�~k$�8�_]�?L����~o�)h�I��}�w��Nb�0�r(���2����P�T�ϒ2�X��.�6��CM��'��@Zp���O"�&�c��Z�5��+i����W��:��1�_�����m&ٶRG�2���P�:=[>h�P4���_3rdY(O��
G��PH��c`�R�LDt`_�uK�g�d�}}���L}B2�fV�e�Ō:�{+�5e#J�t���ɳ��m�n�<F��J��#�c�M����>Uk���������1U�$���%��<=�*�j<���U1��d3y�#�l�D<b�S[n=�%��̘SG�a8�rw�뿁� �Т�dŅ��Z�{�}2�E4=�"u�n����n��s�ڊc��}wr�+��֏�^��8B*�%��k�ވ�5/���A����n�x�-q�4�Ҧ,(p��x��	�N�}���ң�6��?�wC}5x����pq#,L��}�⷏_^���/;�6�6ݽ�I<Kuj��ǒ��LD���@���.~
�_J7��֥�H����c�S�|���~�BR�}��l���%���Y*3q���\�~>&%�V�b^S�?{�t��M��۟~����_o��֫u��t��Aü9�E��k$����Y|o�A��� p���[��F��M?l%ھ�ȵaSQ�!��\v��F��eݝ�
�b�"���]�R�t=y?Q���Z��5���%�e���i�_T'����A˼�����B�i:G��fQ	�L��5*!�=I��H���혐��9�ЭT��wS�^q�����?R�i �4���q�Ԡ^l!�s�\�4&�^�^E6�S�n�d8II�z,RH��Q��̴�wb6��+����PY��J���1�7Pj��	�7���Cz錛��K��/�V����[yg����ݑY���!���K�%mɫ�P���&Â#��7iX0�,��d��^m��,���˺�������qQ��U48��8ujhg�̄������_����Jd���12R���R�i "Sz�|�K��r!���	��ǃ(�a�I^��3)��4��R���јnG�(�iA�f�;H��E��u'Ȇ7�MI�4ZoK���r�0t��!i�ޔ��� �襆	�&)̞q�1��e�k�Mq@/����ݒ	�O���]�>D�4_�bS,�3�T@w3�pMϺ���X�t}QI�PT+٭+�ǯXRl1�΅O���l��G�#ې�AI�.�ǣ����.�����_��VV]�P\�i�$|\쿣(����Fؾ���/�,�XIe��d��h
a�0";�$$#nr�8u6��
T��^��^@Yax�q-5�WɹOnX�_��ҁZ��TXܡDn���ߐ��
tl�I
/�ᦕ�.iC|5�ʗ�b��l���&�5��~�כNj���������F���lp˔E�Ű0�p��n��QU��@^Y�U�z������7�>��?2��H��~{�J���ӫ�����r���|̓��ʗhL��Ť�A����*�-y�"*Q�.��|kP}�����iX���������W��-v��A���+?��K�Ӂ�E�&]qt�MBh�J�\ #(3�Wpe_k:ҏz��2e+��5�:�0&�)�>syN�i3�'���j��-
c��d����~�V��St�r��%g'&8�ށFk����t>�����hl�$�U����l9	��*Q�44��a����<#a���!/V?̿q��%[y6�0����`�G�r���rDҾ!�V�2����]);���?Ζ�1���� ǳ�*�J��/�6a��2i1���nʑ��Z��hU��DS�Z����G�ǯO:��q[|�9y�&e�/Ȏ���+���Q�O-J�������B8�ί+�0��]�zQ'ʁD���V�R�4)@��Ebօ��e�]�|�5�Fԭ���T@O�*��0�v�U��ޣ��	�g�i��TL��-(�W%F.V�Ĉ������[R�T?
��0Mg��E")�ƿ��Sa�2���\͂j����١�+Ղrp�|��Xז�f~�K�����(����V��w7b�=[s�(���[�)��Mο��|���lm�L[Hd`&�y������6N��q�����ͨ=��~<����-�^�	N����I��54�^Q-p���eQ����<�J��mL�Ȩ��6Oޘ�O�JZv�b��	ف �d��܂Lu�����xe	U
l����[��4W%r̵�H����n@�a�U��W�'3�/�+�m�X��*��}�m |V�� H21���Z�I�!����-c�ĥ��<�
�82��=Gr8�_��čb��,����or�~���ю0��=����+�>�Ҁ��n�����n����0�����vg�k7�0�i����Kɑ�<��~�(��/��خ���ctY �Pݺu��R����P�1i����n����*Gڨf�U3�7/��4cl����3{J�19�b�uq
0?ċV��6���	�����O��8�)KYt�pu���Е~���h�+�r}i�M�c�3������T_�^i����2ؘ����X~~{��p��ٗNE�W���k���Z�Ǵlt�Z���V�F���_��l}�{2Ԑ^�&�q?s��co���XTJ+���ȗ�J���s#]��S���b@4zT#��Bj���5\㗂ܺF�>9�H%���r{�M�����QG�Y�U�O�nqs�-��)�O�sl~������:�T\H�����y�H�(ҳ8�q��f2�S��H���3�3� ʫ���O�mJp��'h�:�t�xv.�nʿ��E9*o�}J<���\ϋ�������#���TE���q~r���Y*��T2�Yc�X �=&`qh%���p�g|0x�i�~qA�.�zh���o���Wu��4��1����5Wx�=��@
v���DobS��-!�]�+�8x8Xۥ�	�Xu;<z����:�E����̌��0��Q�fwץ�T+�)���}���x6���#���[�����:�b�揑��tY���q�%��-���87B�E���L��h�D�����n
X�]�0շwL��˙�o��B6q�!�a�z����՞��9�Uh�C��+��z�����ЩP�=����f�%Fp����$���R������7����+E�n��f{OJ��vsW�-4�n�N�}|Q/&ӾI������u�k���k:�=��#8��X���>rh�^���rY�F��f�J�1��?F:e�r׼ji�.餩]�|��jDL�Ejw���W���˂�um�$�2�M��0(���������΀N�R7Oʠ�f��/��.��6W�n����Cy�BNEcj�Z�p	���P� ���?�c-T�]B.����YZy2�3D�6͸��ò4Z#}W�?�]H���A���sy������c���RA9FM���LG�?��n��\���x-�U��0���.���ދMOj�R�9DV^��Qۭ*�vgH�u�oBR�8o�
g�ST�����>�Ȩ;识�U����V���X�����?�� ����4����hpq.��ʓ�Hv�ݖr�������AgȾm�؊Nђ��u�'���T����3R˔��)&���	��:=gB�\'�c���S;�\�:�HQ�R�����*�-�xVO���B]����{�������u-�A�d	֦ɱ6�S�ň͢8�?�%*6O-C�@%Y0rX9]�_�Ԏ��؆Ù}����`�%��>�u�@:gI����3�OϞ��t��������zXA^��`'u}�u�w�?���ʃ����ϳ���..
��A��#��9��e��L�?��橁����M����,��M����y��Yh��&�v}]�Sk9�TK�^��x�*�:�+\>�rH��wR�?�k�n���*��B�9��l�='*��`�|;\�f�~�~@��k�x�#O�V�Hw�����n�Q��0Ƒ���!�g'P,�kU�fC\�L�T�N�(cž��n|_�c	���۟��,��e�S�:�6�6��9�����1�[�G��ٶ��p($�7�v�N�K�gbn��=Y��	�� &�p�eAb�7fEB��_��gvSd�U���>��V�b/��z�!�ĳӍ�M,�1Q63�ς���w�������!̾b��)D��眭���`�Wn[r~���	��caXP��VU��HG���Ŀ/����QX�f>��V]J�{ �\	e%O�RPs0�385�/%�F��?A�L�G�;v�pH��b��Pu�`���3g���i.���!���g<¢��]/�ӹ-ef�~�Sܠ�Y:��d'�z��9[�<���ݴ�b|:�	:8(���sQ�^|cE�K����~)���T_�;|?W�^u��Y�r>�tX��kF}�5S�9z����R7V^��x��Oڔ�h/�]�!��񨷱���Q��ѹLڹG-�e��T��S�x3����;�b�P�Q:].%����9}
�*R-I�ç~&wx.�f���}d��H6B�X��{[��A�g����)�� ��?ul�kCY��7��J���*�E�?~�)�i<�]���N�o���E��Xr�o7z�&Dk:
N��I�6�T�HCb�7L\P��K��g���E���_)H�ٓ_���e��'�f����Ik��S�_����WT�;�et;�Ӯ���� �-��k�4]�_ �zF
ζ�������p��]`5�_�0�i�)"t�H�|1gy8�7U*�6�Y�?� �?��,���0��,�)	���k��1�g�88� h��g�v�U<�-�E���۞C	�ӓ^�~����<#���u��-5,��j�JW�>@���7�GF�Q�R�����j��Ժ�m��d�g�����Mx@�p�4.�z�D�S!��_C2G��a��żv�ִ��/�"Q��b�������a�e���ӟ�i�B�zцg/<Պ_�~�X�[�	*�@O��Շ����^�!��х��N,��I��-�>�+%���W	���?��Xp�7�r�6U�P�Q�5>@�Չ�Hx��W����}�܊
���T<Y|���s/��Z;�"6�D���99rԌ�}X_��]�N_�b����d�bR%�{9��x��Gj�H�F~���=lRH��{�УQ�Tv	s�S�b��M�ӟ�Ir�˰E��O�6�&+)��q�^(�`8��ᩕ��-;�zPK�b�X:�,h�Љ���4>�v� RpHf�����<�s>	2�ߝeC�,ܬ=����Y*�a�L�~y��[����r�Ry|��}D�"M�K2<m1�n[�9(S.P�Z#B��J�j�f�2����p�sOi��1��`� �3�-�EsC�tY�a��7U�B߳5��g�L�4L"%S�#�D�(e��h�j�J!�ʴ�p:��|��TN�ߐ�Яz��ݞBE� �W�1U����F۴�'�\�ٛu��M6S�j�Y���	C�_"���������K^�jf�mH��[A�� ��z��2���O��8�7�BO���F'����ow��-h��ht�Qk��z_��O]�����(��18/c�n8��әGz����G�����޴�V�h^?�K��w�hH���:�����)6yOKT�2=��,�u�"M;��}�j��Bg�S#�1�c3q978���,G����b\��:d�;e��R�׈fN�2h7��0���D���E�����7XNy���%VQ��ޛ:p�Sִ�"]��NE�)#C����P,y�Xve��kU����Ƴ4�Rŵd��;4P��16Ì,��!y-�B��`9��u�Ln���4��m��Cgː�C�C��`��z��H�9�}��1�f�Rb���o��א2g�\��LT�Om��
)M�5���AH���B�|e��!N�.0楝�O.����[��R�aKw1JW�� �W��IYIf�煾_�.J	�[1F5[Ō��)xtk͚>0����q��B��~U<����h�B�shwM�
�q�>����^��k�ܖ�m<:B\VY��e
h?�sw�q����If�k��[�4�W6�����Yz8��V�x'P
��,���l��w��A��DLOى-$��x�t��ڮ�Y��g# �8��E�Pz���礷��ZB�(�š�hEtIn�����vy{v������,�q(�nU���9�x�B�5�{���3$�&��z�ǭ�h	{�Ʃ��6a��������^����,W��rx���]��y3c�}�7O"D����gNFc�TH�mT�ei�Y�?%�g:�T��D��fU�n���{	���I��x��Ԧ�����}�� Y�K)˨nu'��0�(�NL�ܷ���a��^��~�oݒ�q�#�_բ�l�p�W���Z�6Y�yƙ;����SK{G^�䆦��-W���_CS�l��W�G��{)�=���9�8�W2O\ɜ,R��leaf����>cm��H��WbEJN/�'��Q����L.u��cI�M�sؘJ��cd	q�:&�h�o��,�i)jL�#���WF�@�R�^��i��/[,�;��١?�ݳ�v���Y�l�J椽ă�F��ך��<�0 jā>66s�}���R9��e�q��c�g/��C��?��'U�LDR�� t�+j^�_�(�ۂZ���t�Z�١��lb��ƒ��[��H�M�8n	���d�c^��%�z�z�2KV�ʌ�v3��\����h�,���^(7��>���~�Z�������-X�R���q���yi�)��i�ꈣ��s���=��,QC <�������N����d�@88>���? ���Tՠ��~��|�ty�U�;���&eIEOѲ*t�V��d.�:�@ʲ���קE����w�K[_ tM��\�S�獣(
�Rc�G+�%X	�E!���~ ��|�[a�Z��	u7�[�ͬ�.��f����M�SM��?�;�=�0́����Fw��G��B�w���I�.԰����� +L&%��T��3�a�I���tAei���s�w�,]$�'�ѝ�b�+��Ĉ��,���M��e�5�Ҍɫ� j��P��x� ��o.*�F$ŒY�>������T5�X�_k(���ʧ��x���S�1>"��מ��ɭ�8_�\w1*̡����}����y�qfّ�����H��N�9E�᠗+�n�����vC�x�eA�u&���c�)vYq�=���(�Gg�Ӿ��l���EÁ������oM:,3���m	�	d?�pϗ�͖�#d�A��r�-�dUJh� :W����������P$�����@��U)e�C�7�X�dz.���g�d�nE������T�R]��X%0��/f]��m�j�㨴ݰ;g��;����@��8���ws_rc=��yrn?q���{���&,ψ���]��l��ur�VIxV
�n�$�ŁH���`�h<��t!J�j�DV��8uIn.fV�j�AUt��v�4�����l㈦5�������h)S
_h�j��W��ni«1�Έ�5cʫ:}��?Q.�R�uH�^���7�@G�����SLL��E$Z֬ai����F��D�eۈC��T��Q_��|^)`��xZ����&ڜ���["_qV.q�d$K1�7�m6j<�5�������x��/�3�����#q� r���3���㻋e�J�8�x��\�W�����d�HF����b�S�A-7o�.h��s;"l7Η�~V"���c���g���j��)7�O�1}�leg��-L�=�o����#�ٔ8=���-EEF-H�$�0�B.�)��J�b5c�BcF��L��IS���N4RtSI�`e��_�g����Ne��%F�F爴A�2t�٢���+5�3
�N1'���L_M1�nΏz6=���,���X7��kX"t�Vg� ��Z�䟧���0��m;m�s#}�����ｭr6�~��{'��.����D�9�-��X�o�Û�;,���_�m�f�+{}u9AL
��av7��a+̯PK� ��T������̞�a�UViV�(�R�KgD:�!@�C@ElH�^��J(J蠀�H	���K"5@(ϝ��{�����+�̙3s�53���+�ے'���~���y"�~���W��\$ڶ������x��������w�@��d>���C���$��;�PbXjl�t<���0�n��+4>�$�c�^H�6j�ڒ���&;�hS-�F���������%H�2�RQ�i��o{q�['�~�_�>!uG� !r����)-[ljh�rέ^Xo�q�:�g�����Qn;�w`d�1�}|���逵B����G�f{�Ƚ��������}�ɞ��K��'��y��&�6��B�tc׸7�{<7��<V�-������0�I�?�����X����hi#��'�7�`��N{������@~|W��l�r����j)a
"�-�,����9[�����V2��{�����4[� ?0F�'0��z�2���e&��_�݀����ZFG����N~�Br��"�Ux��/.=1QOq>X;Q\�����)�~�y1�_����sf�j��35Ʋ@��\�ʊt�..��&��\����F*���ƥ�u�E�F@���ֈ5�<"��z�3��K���k�����[�@$:�H�-X���Dń�}j��j�2ݾ��Xi���r���˧�Nn[���{qJ'�)�B�R�GX8�4�9OV�o�'�Ç]쩃�n�����eŗ��L%{��x+��MS<��ypݡ{�2�Vq��2~�Mm�q3B���A��v��dz�B��d�U��]( ���Q�wґ����P�/�LV^�;�Qys�_�	��k�1^����6�~��0�W��ajK��(F�z�"|��־�F�$T��-=PA����q��<u��Y�&Cy��Z癆E�qX��3�T�5P��J7��hI�чC�KKlE!�>Ã-/{/�&��5������̼�����~�����ΉW����S��:T<�k��]!�>*�������F��z�9���41��8��x�-�x��!�>�>}S-���{Ve��	Tu���N��G(���H	H�;q����<Df�n����U�Oԥq��yD�������e�4qt6��~>(Q�5�g��!�1�#۷YmL�^	4ۉI����O�������<�s��9J%�����҈]=����\
�S'�፾��~������U���♵�3{����T�/�~�� ��c�z4:�MF�.G�T�ѱ��щ�a]V�R]�+�8 �?v�:�z�R�#?���RC�{P�Xo/IL(���7�4=b��Հ�J3�e���y~���֩~���X�^��3���ޱ����f��o�GH��͏z]!+I�>��jC5{�6:����8�N���	��[�GһXq����=��re�߀�f����$,���e�}xu��U��,����F������P�s��X�̧6���Bb��7	-�GGQ^������$'��Y��n@�IOY0�d�<�d8�XA�W�ko��u������ʲ���[��#��,,�̌Uj{]��=�?D�4��v����L<�����o֚[S�ŧ;�U@j����b�X��P�< ǡ��Fq$�sx��*^v���YM#9k�w�w��o��+3��'�ф�,����	����&鹼�Tc�j<��^>|4DX�CK�)@ȪpuM��Ad�8`��f�����!}�����d1����X��=o�4�n4F>B�Ek��{����@�hHb�^d�	�z�AH<�C��PJ�ݮ��T��C��
����t��zUl�R0O��t�q����<��|4!en3�pJ����d���p|����2O��ń�Rs��k&c,��*iu�Y�(��ա|���څz� d�ΖY����/E������Oa��+�F�j����=�R��OT9z���Z|���7�7Z�?L�Pn�C��T9"g���������M'��c������=�3}���L���+TV*����UF�P��T�*?K����B���	+��{v�����)��^m9jd5u�8,ĸ�-�b��H�t���h��:LF	`�4쒤����	�Ĕ�v����7�'Ƹ�!_:n�;%H���o�l��U��t���}��)'�:bzu�'��;�%�=0�\�~x�;x�ܜ&�����/�l~��G�k�+ո�ܺ�&Ǫ���+��zmz�^(��$oD�=8.�� �-�^�~��Cr�{M���'�ķ((}<�@Z��n6�¥M<||`]��K�>��bx�zPEn]w9�Gby,�^��G}J���)r���"1�|����'�0�2{���2�%K�s���*�i�ٕ��(�}�zd�8��t��>��&�m�g~�~�
նZQ\�#S�F�h��ه$(�ZU��(�#�.��i���W����4Ѻ:wȌ�~,�Y�c^z��c��ő�^���K�7�u�y50��#4�>}VA�v"S#f%����ۅ؎������X�p���Mr9K�ݡ��E'�Ā�C��������(�TI.	�۽��`��5V�JU3}^�~��vY��ZG�\C�">0�9'uJ�;�o4���RFܫ`X��O5&-!/�Q�.y�>5٫�0���2�f;��.[6���U�(G2�� BV1`eYZц�~�����)���F/���h�N��:uNn�sٵ�厠��y�������#��]o_����6���e����1�#/]�����|��ջ�չ4�v���~���P�a��Ѓ&�;Q�w�)[�����O��*B���Qn���`$� ���jtU�ã<�X��Q����k�#��p�y.��w��EEH"�;m�P�k}�0Os����[4E�Ri��3V�#E��=|�����Һ�(g9i����w�p�6-�f���Cd��=�R\���ڳ�0#��NQ#�����p�s�S���o�V�!������U����*_9������b1��$�NQ�@��V	�K�u�����o�y�l$;�e���ϳ�U��ɜj!F	9�V��ݗ��.����D��/�3_��
}8�^P�XN��b �������z�bcޔJ���r~��jhvlW��7cxs�C��u��Z-�r� �����<�R����S[��y��^wD���M�[?P8���s.%��Iw�>��l�W�J���FEsN-RO6��> ��$ؙx�R�*���FU��.�. ��A1vt��.:襇8�`�۔5�T9��t��	cr�C��a�u4�G�+g���W��g��E&7��K��84��V{��;���џ�4�߲�E5ZH��FL�տ:5�$v�f $�EX�{�r���b�6��x�/w#i潋@�.yv��� r��ّ�a_	���`Us�9��������L);_���8.���=���ȠI���v
������hN�!�������g��	�M& .����Ti[ߑ�^�#s0�s��T�+�v���}i�[��/�A1�k�UI�h�QM���2�to�evr-���v/���#���Y��t�_rT7@oV���'�M��(����p3�N���|��
wD�P �1.�2(�=�c�̙�Ŕ�>��зz������J�A��ސoP�bh��Pqb���"����]W�2�ۿ�JT�i�wL�qE�1�����0���SW���Q1��3 ������;�a��ӧR��!?�u���9c}0�����r��7B�����~��Z���N��s]�c9L-���W*�ɵD�@K�Ů�k{Q���W�>G$zAH+̃�_�U�B�RP���v��#?���^S'��:��~�qEM�����E<��)��E�Ԯ�a����.��ħ��Z3W�<v���ǔ/��\ĦZ-\ ��������p��
�G}�ە�u׭��2q����Q����l���}�`����<lڙnA��g��}M�
筷4-�g?�MH��2��Q�.�Q���T�݉�;� T#����`^.��&����͒�*H۩���TC�ia�}�����3�r���L�H]�+`<�*�^G�
�[  �߉l��^�mon+��|�"��ŀ^f�)�7����l1R���7�h0QXC��u���h��zG�-�և��0r�f��˫L5{s*"ε��R�����vy��xB`X��lB.�W���;�~p�>��n����;���zM�WX� ����8F��Hߑ̩������ȒX�Բ�a��+��	6�[hW�t%@�tR��Ə�&v��Ét�	��&��:�,�M���F�� DX�MJ�&���Zۥq,}˱`1�D/��K��E咴�V#��}S;K���i�K9�&�W�1|dJ���q ��O�%�q��L��V��x����Ttq;��f�j�!-2k��*�
�dNr�iP*��Bkk��
n�}WV�b<0 ��
������i��qҿ�B ؒU����#��Ђ��UZ����:�LTg��������V`@�q~J�����X��2#Ӏ;���9o�r&\w��9���u^17h��)
�4ִ4` ~�k,�Z"�U� f�� -�/���{e~����$���T�h��8m��Ɲ�''���2�C�K���A�߬��q讶�����n*e�n��G6P��ʸ�x)F`F�I/�(,���D̠�r��r��~U�+ kX7�Z������EIZ2��W�&ҫr��ן������(�U4V�ֱ��W��̩�O�|��m$�"'� 4+��v�D�4#n��?�l��� W����X�I��;]��kS"2�˸V�E�������l�A$y��Aƛ��v8��Jw(w<���=zt�Ⳟ!�u�v��R�(�"�w��Z��L�xH�c�=�g�� 'o�I�> 0A�a��^��$��-�a�O�f��ծ�Q�G����������l�;�ĖZԾ�i5��y��S�І�9�� ��P)Q�D��cӣДҚ�S؉���sh���4Y�"{�E�Z���5��Ch���γaͭ	i�z9�zS�oX��i�c��H@U}Ҟ6�u}҂&�L�}���à/���Z���iX�P.��R�噵�$�鋁�wgg��7$��;�[���|�/�#?��.�����h�ꄱ4 ��3���,��tc���	�W�WG+��Tyt��{o�9Udo�	�H�E{pB˙R��I�C`i��6���˗2�e_O��9�TJ�P|i��~�a����ѱey��Ch��fI��CS�w�@��C�1[��=.�%�8�=���w|�z%DCcȍԷ���b�O���|t[!*��&^�a�xXw�9Z��[;w����Ŝ��� -�ն_ޜ�1���!�s"�8���hI�wd��a@�Bj���JNSL�;| �K'�_S�3��~T!LL�:�؏�P_�W-�ù���?Uj+�ے���Ǭ?�E^e��+αX�z��س��y
T���v7�K:�?G�=-D�1 ��"o*b>���(!��^��b&��������TV50��&����٥f?5	����P�\��YQ����L��u�VʐH��uX�, q�J�q�������k}�l�-���7;��G��<|�E�Nud7��ܭqX]w)���rj�x]��X�T'��(�F?FD�8ӗ�:��݂p��8�$ }���@��.=��kԚy��[���G�بe%G �I���������dJ��8�Kj�,bd�4E������#{u9Y؄�6N 3Q�Mg��͗�ĥiAY��Wˏr�!S����4y�5�Y�q��t��Yh�4笺�������
uڒzfJ�D��r��<wE���>�+P�۵�.��/j(P�������M�$�KE�W��B*�C��� .�[\p@�������߅w�m7�>Q~��Y�V�.0<&|��CW�TW�Zf�W�'��>�B�%�g� �<)w	�T���nt��>�h�� ;K��KQ�*����}�QQb�7��X�p�^��?��1�>�w7վ��/m�5��S��'����ݲ-��X��n8J˝�ƪ���%���{t0�Q���m ����.<,�� l�Z��4n�YD(��F,�A�z~�V�VKp�5Q��̒��F�M,���6��BV���Pŗ;(1�-:�ȞN��:�����5��Ue��r���aX�׃D��s��c�~0�ۂ���b)� �B�:�O4�ރ�j�{n=���֘��[�!���sl��F����玕�)Դ�y�4d�S���]y��9`/ �k|J\�N�L[�n���]�3QH?[��/����>eV��1E@'N?���DxC	��M�J%�U!g���rk�ݿ�������<�������y�ʹ~�y_^d՜n/'s�*A�<��(��@�ڌ�4��� ��� �O@E�_�Z���[�@hꤴ>��mv@p���y�����1$Y��Z�h;���IP��a��<2zϦ+�u���l���n�KI����7��r�u��;����Wzg��izA��@[i��L�>�桲�bVMу��� &��13ty��� g�A3Ji������H�B0���Ru[����'÷�ty����ĽJ�����/y�e&�GH+�#���*�wI��
��V(�μ0u��a��}N9ҟq�*���zMW��9�����pXIS��u�\�`�5bG�lW{��(��:�=�A�C����tvw�|M��cOi86*�IP_G�H��m|��[��ZA�y<����*M�����v�Թ'A��#~JA'[�P���g�2�h��q\�S����.�@��1d �Jl����#j��c֙�����ĭ�H-t�<SDQ���b��u�]�{FX�񡬫�~��B32,�PD�(3F��t�=b�t�E?�7���PKXq���O���J@����r�y�G����>���"�3'�Yj��>��7��B'�?�N�v? ��_�MF� X�\O=��2������2����ώ���&^^|��8�M������g���{���<��8�l��]��4�cy�dSu��ӮM�#�c�P��M7�S�MC.������ [`p�IB�" |et�'�����\r�؝Iv0d���(����s��K�^e��� nZX�l���k��kd���i\"v�>�1�g��q[�,��)����e�k�z.N��c�^*����q�f���$I� K �a�H��['�}��l��鄅� �-l4^��5\Um�NP����8Q�[�|�]�N��sV:yB�;�u|���x(��]�L�-+�W-�f})��Q�_>WEu!�pŭ^�-2��Q;��g=3�)���L��3RP?o?n���W�uHb#�%�de�����qj�h �!��EŸ�c>�m���Lp
8kQ�ss�7aE̬j�������߉��CH�kO��4��^�'u|��Oz�B�:����qY��{a�^�����,/8d���m�sZ�E��u�ϥb�Ll+k�Pop[]B���g{�fN���b*X�kA�5X��_��>h�o��H�p�eeM���A�3~�7qq�/ӷsg�)��s����g�������t�	�>��9�z��˅�E� �)J
�L� 3}��2U��HV���R�
ș��|M���`�7Z�k�uQ�Mf<�����F"%�I���Vw��)#i��4����0�fn����#CW�������HhG.T�Z�l!���]Q�:KQ4��W��no���DB�i�ʶ�v G	�v��U����s:�tS�L�jۜ�+���������ZT:��k�u�$�"=������ȍ��2,��� 5aYWm�CKJ�xQ���!��`%H0DA3f���:��)P���t%Z�άg}a�\�s��t�W�D�������c��W�Ro1�����o�+T�.��u i��.vc�C-�9����(���z�C$��.��FB�����k��a`�Jx�~ԇ�1�y��A|
�D�����ҋ�EK�D��~`9����'f���%if��9p��T�R����;h`�X���.Z	���
$'0Bw�en� \��������$Y�� ^`���	 ��er\����Ux��V̮1pH�K��i��.Jn�I��K�}�פ%b�Ha���
qB�����	���=���e���P���n����A��Go�glv�+�+~_�Q���c,Ș���>�Ǹ�% ݕ&�S5�����Õ�����I������J�k.���.RkR!1�X�H��~�\��KW������F�BB$`�)��{Β�X:�ꄐ[�����MkI��	�@���J��`�ji@���/޳��$$�4qs.��k����Z�7>�<�K+�:���	�<�٫7��������(��Lˠ�j��6b�ī�m6�[V�H�U��<�I��Mg���+45�.��ӡ�<=�wr�Ɣ�d�K�;Q�{f-~Ӌ]��_~ZxC���d?R��m��rD~��Q�� U�U�2�7Pß�K���
o�:�ܲ�w.����
?I��(��:̧"(
�Z�J`6��Ƅ�Po\�����t��9��G�gT�W�
��b;0��u���@��6CQ���̭_����M�V����	���Ã����gy�#�:K�l�г��do �vH	,NM�ZY�������ޓ4^��7P��	\d>�U��ȶ~'UR L�K���r]B=Q�����%6Lkp���٭"����1����B1��> ��E!�j���~l��'���_L�:V'�w�߯�~�3R��oWw���b���dy���OC��M^w}޵��@%ÿ2߮�:�*E���׶]�+�H���h�(�M���P+x� �u�B�;��/���3?���H�#HI���8&�<�n���������˔��t�Ft����
��ftwp7����֓-��Dݴs2h��%L<C�9�C�+h����_�Z�Ǚ�h�Ub�9|�&�+�"Wn�☍\�;��Ѻ����*ɢ��ב�&�}2k��`�\ؓ�p���	d�I��L��}R���C)t9���-�	�g"�F;
zN3i�PL���/3���(u�����GLzc�#�;wm�>���,ga�����[3�/�7ҶGʎp��Hr�+��H�TL�z����,I6�䷙��*N֨@�8�����~�^�za��*��g��y����٫��	��p)�?�
p�^��-9���j��ͼs��D�'��t���T��u���Nv@V?q�[P������uT��3A�^���NUM��DV�����3�|d����}�TM]�V�gtUi��N=O�a_��eg=�܀vN�5p�a9�b�ؽ�x]n0dn��/�I���xk�g9W�^�J�A4��=������˓8�+r�x��6�M�3+�R8��,����P�u\˵�=�j0����*7J2�B�ܿ�&徫B?�_Nb�>�y$=�rǉ�JkabJ^���l���i>|?a��S�H�q;�P� �b̵
Z��f��ʹc�!��@�9��ș�M��R��I�>��@G���hډ<m�W-A����x�\��w�[��؀�E�/v����ʠ�6{p͉������]��h��OL���D�����K<bۃ_w�o� ��ױX�A�|_�hyž޲R��0�9� ��ѓ��®j��3!{��*q_C4`F�Mv�x���_8��d9y�'��s�s��,�4���Y�QCE=K�c4��C;ٕ�J%������`�/0缠5�-k��~lU��;M9�+i�sc:D-_��1K��:��Y����a(���QYY�胉���9O���E9��6ׂ.���kvw����f�Iwf��8�'%�[v����x���!�`�Vpzy�ZS҂���^$���u7�$3'm��@!#��j�~�;��Ꟈ����;�p���#���m|��ע:XJ��Sg{!�
B1�0�$H��� 2�b�U�Q�u�ө��^E\KN@p��R��܇�G�M��N�Ԏ�l����A�c���)���lI�D����"ő/�DM(O��Q�b(��
�U,�=�_��9��1�6�Y�K��g�i	����#{�-�4�Y��:
�'�M,ib*�./��yQ�E3�ֺ��"������ɻ}�����x8�}gl�j�nnHR�E���#u+�����V��f�(�����VoY�ȕjQFg�}� �s�<X�yp#*���9�ڷ�)O�@̇˱���`~��Z{�:�S\�$cEn����(7C۔�i���״?DSNj^v�H)� t�ċ,�H"�ě�h��JeU���U�k�G��ѻ�q��-x�z�%Y���8��:u�mZ�������v���%(�r�
���Q{/:� ���	9Oj��#�Ở�� mk�sMh��������˧�%Id{�xuz:�������u P� @u�|[�%N��Ƞ��h���.��t�=��1�3`}&�9q!�o.Mw��lZHf=皋�G]�S9����������'�CB��d=c�{�eb�cM�c�=���W�T�KT8!HW��@w1Npi�M�si3�ǷҿvF[H�I�%�n�81�Z-lp��ϝo�7$�_6I��t^\�_t��uկ�Յ�WC������_l��1:�zrx��'�$_V2Ɖǻ�h����+���A(�3����e|`����8�)�����ձ�
��q}�e+��KI씍?_@�"��.A�S *^�qT%��`v�H$w�__��Cp4>)Y[�1z��<����v+�1��TwŽ����1`[�k�TT��{�Kz�=1J��ޟ_@�[�:Sɑ��uI�T�Ro����Y�������ނ6�;`�
K������y=�m�]�Xp���B������@UG �ĵZ�&�ڬ*� ���J����6�󛓻nSM�&$&Y%M�[y�}j���<��f���\���D���<8��B�si�F	��|w�=4�$�U|�������8���d<@�_���n2,�J�R��U1�nod	�[���E9��F��`�\�F>���QV�E����P�K��2�ךmt���}�@�N���	(xQ*=P~�u��{?����s �B�um{�����Eo	�b)3e�&Z�7���c�'�QD{����'i���mΟx�����GoJ6��g,ZvҠ%|g�*?5���L��E�fW5�����_�g����?jp�̑���/��\+Tc6ԁ�?#O��@d��h���w�cв~��(���gil����S@�}�@z�R�6�{P�T@�g�tg3V����*��o�$�/_���v��,��~�ʭ�j�eY4�q�����.p�&.��N+�(�i�Z��ɵ뽇��ӱ����w�����Y�|�� �	1ʿ���6c-��"@��(�Y)��1QH��3�ɒ�J��4�@�ˊ<Q�	�#YnS�ލK�בv�.�;��kڋ]�c����F�0G��~~Y%Ij�����|��8fm�����U�U%1Ě��_:�>������e{��)�1��ۈ��l9 ��V��?����Y�����Y������h�� ��g-h�
I_M���Af*���z�^޽sÉ��G	m؀��IM���Z��쓨"XCcttn�Qu_I�r��K�::E!�n�9���>�a�
,>c�����wnlS��j>�t�E��R���X�N��Q c����C�|������8�e���+�jlb�jm�i)G?�a���"����Q�+��hjL���*_�K�$vF�K�L��@ͻ���?�v��e�Tl�n-����������ip�fP���F$�w���Ā\�?Ɉ+e*@3E���K��L�����Ui;���x�V����h��R%v�����VLL�@����y�Z�91���*�؈ن߰�|����9 �a=E�;�nG)� ����
7�
���_~$�7z^r{�b�P��X�=x��)�P�_��b����	�m�Th�ϵe�Ƅ�(���>�y�l�����y�ߢ>#
�n������jsI7����⭶P��X�o7a�NJb����B�ܟ&>/ǰ�����)�U���j�Ij���&��ct¼Iz�k҆|H�@��N���޴jv�o����S����� ��W%wxT)"M�[��h(��C1�9�~��QZk}g�}"�^'+/S��kbn��tSi�jLs~�:)G��ګ�;'{���k���n:��̴���$������sD�32V�d�oU��$�o�l&s�[��1�..��o�{����s_x��n!-p��d��W�ͳ��ފ^a�թ�&U�}��M뎇G*�Y#	Tb��;,�ڿ�ϻ\�>� �� x]h,L����Ag_��]-���5��a���/��n]<�A_�'�t����`L�c��|�K�����5}?>������z��(���������X�r�h�A�en:N�+�����Û�_*qQg��";E��m|i$�S�0J[��7_�ۄ7��.�?�l��%��)˕�PX��)�<���	��S�����I7j9�R����=�m��Xj���N1�^��K�x��3��9o��j�H.���:�d�>�v�lҽ^�-��j�ݹq3k�Ok�~���������0�y����jˆ���ζ�[��N�<�d�J��[����cAA���npk�AD�M	�W�R!���(��R���2���*�t����hK�)�ܮ�B�_�Z����ߴ�;�����C��.�u�rbf��y)	�9�bא%�.{h��n:~�~�Zp�ALg��6{�x=w�K]5���@BN���5%�iÜn��/�dN����>����z��^i2u��0�gb�c��r�c!�UöQ�W�6=W���v�`=�B.�o��ow���q2z��X̴w�{�Z�c5!��y-t����*�\hU\s���AIo2�Kk��_��OTu,�RttP �b��h쵛w�t�������0n-����"��l��s�I�?pW��*^ĳh��k�[���J#L.\��H��E~ގ�aj�1x�'�<�+�}������p�Ixn3}B�����$S~߂�2$��_^ɾ�#�I�E��z]ŗI6&�]�[T�Nb����y	�Iy�"��NPTT����ъ�t~�F?5y���X}�)��;l�JX'#ކ��o�тs=�;�e�D�7��UG��J�)�STUϾ�=��Й��p�Z�tդ���ݯ��R�?�w��FxF�Џ� �}kf��Z�4&���Ղ�}�T�D��2��{�^$�b�M��9�m�	��AI�Z֓ۮ=~�:�0ӱM�1���E�)r����Ia��P��� qsm�
G5�˗ώ��zę�V�*�;t�h�
n`޲���u��χ�SV����.|b�Bk�ϫ �b(N���GY�8���_em��� ��1��%���+�^$��l������'���Fꂲ���A��E���w��]�r��j �b���պ6;���1U���,0@�1)Q��9tl>m���ѳf܎�g�B�&\���������ʶ��� �Mr1�A'�r���Z�����I�]L��%���?�H�s��J���'��	s%���bd�<�$zec����#c9�Q)[L4C2�#k���%D���U�u!�}w�J�o�g�m� v1DW��V�>�2��&	i���s7�����U�̈������:�lY�c阊�=�Џ�8h���l�s!��GG*���o�FOqQ���?2�x�B�4#���]gY��7|��7����K�v3農���B������g�M�Ea��%���i�_����V���8�)�2_��#� ��ƥI��D�1�W��}e᫧:���_��hp�RD��a���@�|�M��S\���m[��@�u	��
�`��)�M_x�W�s^����D�*_:\��8(��y�oC)^}��eͷ�Q��i�޾ZHcDWK�A	@N��-��L�"�N���wr$�>~�������D�."�N?��!��<���
�����:��L��x"o�:��f鄇h)=� ʚ �[��݅�@���R�	Q�>%��#~~�{r�� ;8d��戀��q�w�������
Y� W�}-�}��XZ�QS��5z
d�M!7��'}Z��\� �lT����ga6u>+������������O���s�VcXYPn��s)6.�����ut�o������mV�<{F��z�ա_ �ګ�,�S�qQ����x�5�Pn��K�4]��@�K���.�)k���v�cJ�Y��-}�s���V�Z}N�]����h��b���,���~׾(��v@v��R�sXR��V~�r\��W7[���"wn��ʰ ����?W45����b�� ��ٗ��Z�N�փ��-�/��n~�.=��Jox��3��ɔ��3�wҹ��(% ��++&	(تr�t��]��?���n�����7��)3(v�s�Vc�`�z��qq����f�á��jy���Iw_��;�4�8YX�ה�Z�(?5���C���>{F��?��^AK������Tr��s�9,�����Ɯ�3(�%���37�Ş�4�ݓ[U���#�0�e�w��gcaYC�݌g.�=:��2�(��H����7���p��-���4\!���xk3��M]���/&J�b{zj	{����5��w����י����2{8��]Tp�n�q��ʋB�p[�{���9�����_���|�6RRي��8N]o��\�.�N\MJ�v�H�ON�֫~{�3�?�$�L�:a��>��Kg�;�xx��gKFB�t���?<\!y�>�f�[Վ���y��]�>�
Ƨx�ι��}{�оj[�f
g������S<�{x�)��(k��?cM@��#��%]��7jD�9J�y�@.��k�م�Bm]������F�]�^�T�2.���IBy�7���R�u�q5?n	yU9-cWS��zII��0K{��'���'��n5���*���ollM0Y3�<t����!4
�.����F�oK�G��.<̪���/?D_J�7�X5ʫ��v�>���E��S�'y�ؔ�j<��:����Gl�?f��.�m���}���z�����:�o��,1,M�n%4����.���KL"귶E�v_A\G8i[���r�D�W涺ԅ�GF輸�="z�:��d=���������aGBX����
^ʷ���&?���r�5���8>�_C�i_����?�"�|���z�v��"���Ԛ��3���P�߻JV�{�s|�gU�ľ�[���p!#�c�N�z�TH�v��1���pm9H�v�B����AJ��#�w�,YzD�r��K����Z����Jb'ٽa���-r_�o�~<��`SP»���-�p����x'>�ɲ�E�E33潊��rΨ(�ƭ'3��A��lW��C���X��ٵiji�����H�[�Ė��Jaۺ�?�>WX앞�w�l��Z��D�T�<-�_�*V!�i	Jmv��m���j��t�u���C�_nT���'Y��mM�ꉂ��g����>-����Zפ�x���_�,�O��H��|�o{/�b����L[���_��<"�l��'?�˾�j�\M,�IQ�s��s��~�Ob��U<�M2���A4~�G�Pa���#W��F�ޅ���w�%�����%E�ƅ��������x���p���Sȍ"������m��C��x��4g�l������ϛՈ��t�oWGc��#�q:�D|v7����#�"�voI�Ռ3�;�b��lz�N�\ˇ�/�O{���ń5̣̜�����mf|�!�Ac��=jtB��>��j��h��־܆s���y���KT�R��q��MfW;�M�m!�T0�Z43:�V^�^aQ=ȦT����8we�O�<�e\<��(����}��5����|����u�gK�%��E�=(R�Ԛ���bW9�}-���6��VZ��Yb��g�k�с��G^�ֱo9]g��S<��H��~��j����h�3)ɫ����@(TM�	��Z Xa��"a�_B�����@|Sb�.Ņ)�6~m���w(.�m�X1uxL����A���џĐ2�G�FZW��?�O|�7	�F��?�U�&]>�sv�m+H���I8X�w���?�FtGe|�}�b�/�����F��_<�3lZ��*�/�E����r��<�Ɛ���K����у�=���D��6��9��o��v����j�Y��cU*�)�oz����ډR-yE�f+��3�zi(��X��_��3��ok�&?��lY3�=�Nd6�t�L�4��޽M��E�I�?��Αз�J����ixX��{�����z��$�6R���[�4������S T���Ӵ���KU�%��Ψ�W�M�Tx	,�� ��d�e~}i�8M��(�O�P���hG�	�1�d������{�$���F���u������7�)�1�ѓ12�E�=j�l��vzq���>*�u=�?�%Qf�OL�lם�c�<@���?�]�����<���l�RG^H���v4��t��3-vj���tq�n~dM�xh��ɮ.���pj1���Vt+c��L�4G:���sc�k�+{����j����XQ����8�-Gl���m$��8��l���v|eʝ�����͕���:��#�f]@��A�v�+	�}$(E}S�=-9A���66���۞�7;�20�W^%�	m��5g����t�������?��l�o�(IGw��I����P��gr�9d�o`2�'�7r�c��>��-]�P·���^c_`_PA(=��]���c��:$��͛6"�YE$|�ͼ���!gb��׹$JX�IND��1�u�!�?��r=���7���5�+q�q�s��[{۰��g:��{�A87����Iv;n8u�՛��uϓ�_�M���>(j��h���GzsPo�fl���A�Z	
��ƩT����������ݽ����o��z��?���P	݄�N�R���q�pJ�ZH5�r�Ƙ:��D19��\Ɲq)Br�}3B��m�����9��k������}�?>�����y��콟�_{?ϳ�VLٝ����*.P�;0ݏ�:.����FO'��H��Da���`F֩���͟�u�\��I�J���,ª����&��o�t�4���d��U:�����:�[W��7�ݲ'�����ډƇ��i;�;>&5e�C�'�'��zm
���F�k,�Xg&H{�\�C�~}����'�Y�/�
5�I:���c�'�Iϩ]nM:�i���h�$��@pAn]D;_˳!'�O�l)o�LUG˓��RU���ߚ���"�Sfg��y_@UJ���h��NgE��/�������'��E��gwr�����x\���)z�5P�'ڢ���y3V04���.����dX�]�h�[>k�컵G�p_����Lf��yJt���Zϯ?�4F8@__�z�?�vK/�`���^�8��y�A�/��o[M�%�(��Z5sp�����8I��_�2&C�����2��G�h
ޅ�s�g��]���ۍ��>���Ά��ϕ�� ��]5E��� b���&��������a�|�̳�����CPt�E�J���8g�޲��:���d��u¥�@ae_�Ul�ǯ$[��?�����\����}��t���F�ڌ��O���ࣇi2�"NǨ���UA�	�Llqcf�v���#��NЪ"���+�n�<%ҫ�׹Y��g����y'�e5�>��^uv��YoO�h�&���9���{�c�Ǚ&���\�oY7.�\p7��[���)���m�������7��Q�98��V�ŗh77�^�3��um�����g������Y�^p*�mK
���	@`�~�}�EX��~��>O�+}�Y���IbA
D��2s2�������o2O�y>K�P�`��B��yv��EJ����[ ����%C.�����h�^����0Z!k�CL��I�ͤ��F=	f����_���cw�4S�\���'���Tz�'��'�0�՚G�ӿU7�o~� �FS��^t���X)7c�(� ��U���k��,�[�Ӥ�+= ���`�F�דB+���D��t�v�?���|@�ƓPG|2���Փ~��SƊ)&���{[7�"�@˴8�(�c�d���O怈�g�����q@�M��O�Y)>j�h��H~T�>ɲ艕���"a+%p>�7�T�fr���QRt<�Cz��z��{��w��o���~s�K���ۊR@����wΒ�4�[�����S5�˳��5b��i���/�O2��^|������Tx~T��Fd���_��-W8���z�u]�Q���|K����I��hY�
ώ_n5�~O�T8[8�P��~z%�T�	n*����� B��B,����`�f[[2く$ō�hy�������c�j��)9�����09� �š6���p1��,�1��ͼ�m�/��^�nlf8h}�������V��t��&n��~�|ŉ(�ɪS��Hg���xxc��s!uN���=�ƎE�v|�}�9����%o��?L����ݦ���_�s���!�{O;���..������ڜ͵��7�z�:P����9��=��=-��'� �jՃڳ��9Okt���aߌ���o�l���VJ��������v&q�*�|1�χ�o����~Cm��L���"F���JF@N�e�1ӑI>x�ox��s��������hw���{i������K~_7�7���k�δ����&���|!S�Rq���\�|��,а���*l���ϵ늏	�K$���*>�9F�5��>�0_�G2�/���G\��ʳ�>���Zڕ�X����L�Gd���H������I��N���;���*ߖvfpW|��4s��������܇٥>�أܸ�������<瞄�ŮN���m l7�6�������J=�_qk���"���a�ƧCS��L��~���)���V��ǡ�M)K7���uk�~�>��큨����^����qt'}xTK��usa\H�Ю��J}Ŷ2!N���`C�R��(d���hE�?��՟!a��q�#A��[�K"��7��;��� G��UT20$t�wxR��}�r�r�s��m2�t���i��0k=�px�ϟ{�)v뙗/����s�(���K�C������1q���e5_��O��}n'�x�o�X�����<�t=LD"X(����Z���K�O�½�i[��g�>��$_�&�>��l�a��%���. r,�b��2����k������l���}�����ot�vvޣOyf�w6l��a���Yh��"�M>M9�_�P[8�Ԧ�DȬ`<�=R��a���x�+ ,�7R5���fT}���#�xy�;���cJ6G�M� �D��u��'&�/�,�����QR�L��'DP��n��D�ٚ���|�y[k xW�l�����X+!m���(��i ���ތq�M��hG���zN2�Iwj6��x����Ĉ�?z٩�g��˅��?-�SދAH�5�l� B�3�1�����3�k�1NF�Ue�.H��L	ءj�\�X- �ۏn�p�yߵ��n;��#��������������4�8����U��YӳG�d�,'����A\���Gt-��x[|��R��H�����﵏0����/�v5���9���P�E9�����P�>��X����@b��^}�c��IC�ӈ�$����������+���<�F΃�+[72��l�0��
\�a+)�ux��e�m1��ƺ�u�h�[��L�Y�XM��������ӗ��3��k�Z0f���C@!`�S*�A+����Z7�g��,�3'�ioUS*��6/.����؋�>	��}��f�K[I��?�"�ɍ��a<~��ļ疵`_1 ؆�U�4�n��)E�iuA3��$=�+6œ_�B9�#C[�8�2Iغ�wC��ĹsN������nss�P��=�X�@�A`X���S�i��'g��{_�Bj�UB'w�ί���]� @4?�zB������/�R}\�A}5Ҙj��o�X����l��%7��{BwpL��m��|�u��r�6&�b����`�UL�Y��_����,PnL],���L�$4��$�o�W=�9e�_,-�?PԀļ���WuR>�V�� AD�Y�nA���P�X��ԟt)��Z���i�4�DJ����b�ߐi��^}b�Wǅi�a�����҄I�M�"��>����R��<�(w;����	w>;��5�w����eeV��D�����{�d��e+T,h�$�	�:{#n�6IKK�)����B4��5����5tjQ�@>oz��}6�$�RxM,w#�5(?ϟ�F,�r�Mq%-\B���>��s�wFNB��40�չ'這�Q`�L�� ��љL��C�V�
dV��BZu^�Y�u}�O�KY�WCrZӆ�o�]a�''�o�;�U��Wjv�:W;t�g�Vl��FEn����ԴND�Ű�<�[��S�g�kX�X�)�n�ԛ"�+k�^��9O�..+P�f~���s)��ؓF'C�`��}��(��6*%�������u�t�O4��t������ɚZ�JZ�[�7��U<�E��Ĺ%!���f���G��PEfN+�PI1��� ��4:BҀ#l��(��$�cf���5a^�!-�B3�c�|���{��ú�F��ʗ3+G
���6C�!�tZO���#��+���Å�BZ�<��5:�Ҭ�75�|��� 7��C,�!ۤ ��҂'G�#���<*��d#���A��.���%��#R�
<h�l�ş/�ѸXo��}!��xmh山�~?f������j	�K���T���L*N�Y�%��0�k�'\�|2+���h��3���ڢ)��Y���O�G���˚�WlZO�8>_��j��~Ya�ƶ��_zA��yV�;�����[s���;��{����V�j��g=)��Q3�FJ`%a��T�G�kV���Ԁj�H���� �5/��DljW�}���(���%2,l�	jω�Z2U�iB{���j�$T���wz�F�a�#^j�Z\�8P�w+��Щ��Ǭ�=�����}��mJx�{��O$7��ܨ9�bpPF���X����f��{��O=z���l t�n�X�MǨ���кɯW�9.t9_���"��B��ǫ!��n���9n@GT\1tm�����i7���V�D�nB��Ʌ4��G���H��\�
-�3׌<�-�.�DӪr�����SI�������)��^+�����,4�{��f�~@\;6г�"'_l�v�#�
ǫ��`��DO�z���;"����SRܢ�
�rm�w+�_E}$��yl�~����ۀ�����tsV'�w!#17N��j*L��oK���"|q-��{��>�>KԶ[Lc�����S�T�]��R������˚ׯ�`F���dq�����JB�>�D�)B��:��4����!�c$DǓa�(� �ɳ/W$V-w|ծ���YRL���]�矾Q:R���bU�7%�L�+�WO�
��Q(o�R�Q99�~��q�Ҹg7�CZA��Po���)��v}y���Z�rO�)"H���+T7��V�Mm�����˰(�>�+�`R��o}"&�[pK=�Ӆ�^i���L�d��0Aǟfe�3w�:K=�-�d��I�[��e��E6!!��sH�kT�%��� �5fz@�P�*Z�8�<V"�A��Ʌ�6E��y��\��KlZ��$�:>��R��a�nn������Zz���7��i��X?ہ�� ��d�!��`gٜ��ѭ�Z3����(��>������q-�A�H����%r\ͫ`|�^-Ά�{�&T�_h�9:FS�Ѭ2�(�G�C�mW�\��c�����f�a�CT�%���U̬[,������Bl��R/SV��]`[� im��]�>s�Y�%�]S0��R�u�kOKG^���(�Y3U^؊��M	@Ϊz��"��~�ȧ߹{W�ۘ���Lor��!)�=��c�F��ӧ��iXx��͔���a���ѐ�N�}c+��b/� G���� ����`{V��2�|U �=�Ɨ#�6Y��u�2��~�)`���{���/�߁~w�7�r^��4V�E=��_�%>p�YX���?�c��� ��>0������u��}��3E�w���afE�z���kR��_��?���C(��l{���S_������mւ��unF˧�O���u%��v� �.`F��� DM���^�%���鋺CĕJt�h��{�lQ�SW>��Ea>*)�����c�==��}2�����|���as���3�tm���aBF-ͫ�xh�F3��b���^���ga�HXt�~�p�6}��9_�#�g��ܵ*%R�˘B��R����ܓ�(�b�"�Hd$�-����@�:��u�jJ\�����|�F2X1g�3W�}�2�HV�;|��9B�p�c�I�TjO��f��Q�7A.����K��~]U�=C(�z�M�R���y��y*�	���\Yq�l
X64�3��!���O��q����琚�W��g|j=Vuz�%�؇��,�����҃�3����L��]�G��3���O��T
��e�y�ȴ��.,ww�u	�<�y��	v3��ɯ�:Oɻ�T��t�dV唴����罋��u�dn��,a�i��ʩ�Bx��e[�b���)�;�RU��*_�GP���Щ�wa����>�Y[l��`LF�ɂ���Cuم���l��k]�S����0��#ֿ���3����)�����T��1cp��Bi�sv�r�?:��Y��������:���!2�j�Z�u���@��/�I�i� �«�4]��f؜�F����Z���U�u���ԃ��o��'��3�<n8�X}l6Џ'�����_t�r����ċ�OXz��_��M�^�׏�su�{�7v+�G��(bkk{Ğ�|���%�7l�~�=0���{Vvʜ��� �����J��y��^?����zd��0&�o�`o�s��TϞ�U�����b@��N��Tw��n�MJr_��.����M����u�<���f|��v <
j�*v�S�޿C�K�4�q\�:�8���Tk�K��{��}.��Z�)B��wq�F0��Yr|�c�]����
X3���gW�m������<(�[��E�h"Ǒ�{�^Y�x��V�W����}��<6�F�C�x�"{�i�	Nj���.�B��J��4�����҃�е`
�2�!��xSWd��^�e�6�J��>�,B�^���8�'M6F'f�5%%� ��{���[�o��#+��؇��rət��,���ڑ��+�'fĖ��6�N��q6@�����"EIOz.��,ao�b@��q��{�4R�~�?5��4�,f52[i�+	���z������Dƫ���\�}X�P|��EAa�OH{�P[/�%�	y�$ ����&�!E.̍^�ڡ뢑|!j�VN��YF�U��}��s���\\5H����Im��I7�SS��>����Y��&H4n��-���n��Z`2}����%��κ���vɁ
���1۩X��v>M�rt�H�w���n�7	C0W�h����X�ʑ�{����t��3��?�������"���s-(B�w^�<��vt�S%<4�0]}h��D���M�X����|ĵ�&�T��h���_�%k�������l��I��0����=i.���\��s���`���%ȷ�����$`Z6�TU��"�X�F�V�m���i�|�F�A/\N�&
:�`��TJ�}� �}T��Cb>ח"T���&ȌY�ݳ�z��c��^���D���]�ri�ң#& ���Gh����se��7lN��Z����vJ��s�Ņ� ��Qo�x� ����e64t��S� )z����Vn@z0��M�,D$M��{�������ޥ��1���X(v�ц���#���^�۾�%Rb)a�:��WV%��mY�����-)4JA%� 0��A5y�7����\V�8�)>u��(^����v��W���"���@jV<eb�>ء:�Hzj���`��j7�F���f���1�E-�W���U�E�1ʾ6���Y�>[�}�E}�8i)�S
3��^fq2EØ�`�8��pA@�n&���}|դnw+e�V��J�>�}�������Y!1-9�s�& ��Z�������q҂.���+�\|߉��41���>��؇}7y�,�/D��-�D�5�f�Dqx���9��Q�� �&FNZ�����`�u߿eG(�X�r���a(��l<�����F)�V��G�|���ZJF�%v�-܁��қ0Nf��E�C�U7����k�)���.�	���g��z���+;$�k);ʁ��^��!�S���1jb9)��)�>bJj��
�grD�����Oos�Xo��G��i�:��W�����6z�73�jx3����>�?�e-A�C7B ���b�7���J���i��\$J`,����R��k; ���Y���S ��s�K�E*hҳ�@�\?��V/|�uQ>�x���{#<�8"�1[}U�E�`$N��E�� �g�@�{1_��z�/�]�� ��"��i/뇇+9����,�}�*����R��M��e�a��c��5��Z�
���'❵�Uv��n�ӕ�A�¨(��m;�Y�0�_Kz�ѓ�F[Q��:Q��#(gzx|��!{Q+���=���yxo/0w//1�▎Z?4z�������'���dqi!��D*���mr�:�ܴ�wD���&&���k��WoK���r����63�E��,R��rn���c��͝	�=dN3#!&�n�@W����b�����>�+��S<�,;�]���^�]�Hm ��r#�	[C���3ZJ�	>�}�������$_o��jh��[P���I2�
�4����_f�ZG�o-��g��Z"!��^+����c(���^�R��ǣ���9i���]i��[1~���'����]�߆�g���7�	������}�l�qm�'8U4�Gk�~]��'YA����5��e�.ktz�\��!$�U��o�Ё���'��81��]���g�ֈ��J�^���C���$EkT#�k ���a�������l�-���T��Q@�Ĩf8�em'�u��~���W�S��)�; o���S�̛�����1$|]�����`����f��=�y>T"v����4%�	��_�2o�e��bz���8(��I��v�ˍ�}�/��W���G\ ��D�yR��L�����m}��Yk������l`qT�_�(�����4g�'�c5��$j,��(:�e��CN���ڏ9W4S��e�?&(=|>;�d����N�	��%��oQ��){\,�V��8���o�:˂��8����]�q�T~n�|W�"�D��M1�l�!s�Ă��'&�ɛ����E�r��9�F�e����:^]i]�a$��@��;�yM���dh@� `�m�x]*�X���:�q����o��K��U�R
j��S*���4���5����]��oUi��;�»��	����x@�Z��y`L;��4��t�A%qT��b�����D�j�t�"�s�L�!��1}4a����`6����ں�n��\D��j��I}��qك�[�u'ʍyC���S �^!`�^��v�_�Ms��N�%Rx�U3��}���{%�(�d^�ӏ��ij��7�RS�X[�b��U���m�P_
���������*�[����*\T�<X�3 �I�*���9uX;`y+ሄz=��I���;�{N��H����|ח����|��u�d��G �t�'��T;$E�b��D=���8�	��+Y'�&�e�� ��9qq�e���	f	���`���gR�s][lr�����f/��g �F�z�� ��a��K���0�P'��~샧�Kn�X��w�̙i��Y��S��>|����v h����*� ئ'tPE�?�wݙD�������WM��-"�[��x�s�p��]�������ѯz�}Q��;���Q��	��=�ܓ��B�k<����rg�fҽoT^�����o�^� �l\���2�U��i{�g��R��.�=9F����#�e�R�Mˑ�T����/1���8����y��3�E!�ߴ�Ij���uj��h'5�%�GCh��}<��HT�y�� "6��v;`�Mno��L�N�8�W�#3f��<"����$>���W��*36�g`���i=���s������
��;�}��p�d~���>���/�X�ґ�#�Y�9෥��H��W�۷\7zntspEK�D�-�)��y�F�v ����j��Sƴ�X�76�HW�e�������\�G����v���7��7m�����n#_�\ch��D� �(6ࡏD�e=4����	��3w܆4��3~>yl���F�3�9���&?ieluh]g}���`F5�[ۛ��(��ۀ�����f#<N;Ǡ�d�*@�a��Շc�Ѳ�_�� �B�;��%�~uVr���?w����"!O�u����u�>ƋH���;̶d��q���s��6��7����2F7G����>����G���3��TQ}V��1H{EP0�����n�[b��(�::���v�F�@~�){�X8��g�A������04V�5q�:��ow�\�Mֻ]��I)"��:ڤ`��C�D��8�ʛҜ�R�����5ЈQH̰�޼3��K�Kqr;�^�0�0S������k��<�q��R�K���s'-�NA�S����5�þ�7�3��K��ݤ�X�t��Ge_�J4P���U}���jFʣ��G�ň}��:��v�%[�Ja#0W�"^�*����7�a]Κ�Κ#�\�F%/?��MΥ�����=A���:o	��<:-�����ژ���Gci2��`\�|ձ�'�{�D���Gy_b=[�d.����VD����B�А4����������1P��a�r�S�a�`[�Pp#!�Գx�Y�~�$K��3����-��̓�Ԩ��H�� }��Dzwb��m>�O�/��X�q�X���A�/�t$�f����ai��jC
�|�����2���(����u���;���v,��JY{m��.��|b���4W�z����}PaS|����A{9���Hj�9S=��d���xܰ˸�ĘZ-%�A�L�~�86���ߗ Z:�au�5�w����m�tC<݂���v�p5�v�dp�*��X��C�1�TQ��v����'�.����������o����E!���Щ�N��3��D<ץz#7�����6�Br��yi m�w�MM)q�5�y�H1��l�����Lp�����T�A���:��+�eG51H�?'��Uu6_���8�/��X��9�t�`�Snա��	�XR᪏4m������� �=!��F�*�Z�6�<��Q��������,r]���r��52��߄�J8�G���=�$MDѹ^8�������� �:�aX�My|����z���
ER�]���W
��p?���o|_�����k��:*+h�OJ2움���*�@�m�{�~��+�Ƭ��D��PT˸/٘s����\6���^N�2%)�.�q�XRv��Q&:���?�Q��DZኋ����}���_E�|V�^����?��E��[ p)�y��;��d�*MØ�1�n�؞�����v�ϙ��4��qJ�ӻT�sp��|4��J��	���V�fn�H\.҃��jg��_\|�$��?�rں�0�m?/a����}��^��h�ƿ(��t���k�志� �I��']�J4H���;�����jo��ŗ��'�-�]7MU�Xz#LD��]����mZ}�1�!S�J/¾�`��{� �[m�?th\��� �ɣz��=���}3�]�_z?6GR���f�'l�U���������k��7����Пa�
���[�A�V���ǉS���#�A��n <_�0n:JT���q�I4�+�Xd+��i�.�xa��2H�BQޓ�X#}a],�����]��=#d�uo-kݸ��vK<��$�j�oi����xs�6�=MbQ4l0"��k??��x{��8)�H��C��W_E�n��%���{!��/o��I�w�{��p!���&>53��>фk1G���,��i'��7�6\4T|�z@���\Mx��&F�'N�w��ðBb˗���h+Iɽ�Kwţ�<�C��׋ݒ��eA L�^zw�T\�܆�ҟ�|���˫>^�P��\{z���8d&.��nMP��������(d�����	���!O�\� HEU �w�/�ﲯ�1c��P�}͞���CQ`���!D����1=���\{㑴e�������p�hq&I��0�}�� �5��J�eL����k�Y�2a� מ��bΨ	ݪ�_)?j5�;c��L�]̪�`o�I_�m`H��b���	����1*r*��j�[ťh��V",S:ڶ
N��*�݌k��V�HDJ%���胦���H�sg}җ�˔)�:/�}�ʦ
K�ݓ����e�U,�Q�H����Ef���x�gJ� 'e٩��<���jЃ]�������`įu�o����n�����3E{D�*S4o�������Z�٣	��r��}��	�Aفm�P�\�y������YK�,�x�]%* `�tg���t�����X�¨�5��(}2O�^Sai�Z �dيJ"��8���"{QZP����0���2�R˜?G����e#Y�8U�m�:��s��_}~�Ud�'54�^ ٮ�L����S�&N��2��\�����ŷ��c�.���f^cƷ��)�Hs��M���$�z�h�y��M7C�E��qR�<
�q#IƝ1={�`s��7�],p%3���4��v{{�,�r�'��M�'�	'.���F�+H�к6�a؊�pA��Y�ڵ�3U���>�o���1M�w�G�{��ٶ��Z����:���W�e��~�J4j�'�Flέ*ܕ��U�\vE��*���U��n��g���S���½��ى'$q��|xF�ڹ�:�J��f�VuEF���w/�Wĵ��h{�J��WK�4��Mpu8����g%&��$��vfA��M�1վ��	��O��_�`��&&G�F�*FH�$	��|����H�x���>l��ths�1�E�W��4r.�S�E�CH4�@ܩ�GG__ �
��"!�ta���Ǵg�ܶ8�D���˗�V�L�卋���$��,�-:��0>��0$W����eCܫ�io�z�9d|�m����hCJ���B��L���	�P,�_��.Bs���t��kĩ{T��8#*������۰�ZZ�6@���l<�WѠ���Ky����p��}�8�X����~E����"ި�<�y�V�_r)a��zU���bo��4Wb���`CS�=���3=t�KZ��;����n%����W{�n�C���ӹ�2�UA�կw��R�N.i`�������֣Ao˽�߷}��Jl�Ԑ��Xh�p�7�ё�lK$u$Xu-���ϖ�@�>�):C����B�m�C#��,��ՆJ���x�i�HE矛���� G�9G	�&1���#���ݼ��Ǎk,bP�[1_���C_A22�n����ry�e_i�!�e�}N�d��
4G`}�"}���J��������6��mR�Y�m���/�Z���àU�h�rgGY�* �j;m���їL����Yg��*ۡ��-&W��D�\��!N�}�U��s�� 7�h��o����@f�ZC�6\�.�w�h�o����&�4§�W��v��##��
Y�c0t���Z �Ԕ�i%E��PgE@�m�ކ������s�O�⢉��u����O�v�؜k��<���j��:ۉ!���]�����!�F�Zs�L�gW����d��q�BJ���Z>�<-�!����0L��0���b�۪�Z/B�%��|�O������>`�� \�����76�喫'm����������K��y�g�@wF���R�)t�^�5�S�TO	U ���a��Y�m7��R^;-�Ь���T	�Q����zH�Dq��B�]Hc^�"l��f�O�^�Z)�cya�G{¸��B��u�Ĵ���?1�ϑ^	���,2V�C���n� ��.���Mz��sj��=�8���P9sꋾZ���}=�U�q7���%���O�c� �c0�=R{ч����m6t`5���>����:�����u�P���I�2��*�����N�b=����H��v���~rɋpibǗe�v�i�r��Z���b���0�� �yqV�݁S�d�r,d��1m���҄{9ֵ�DZ(���R2�,|\��ڒsc�=�V���dO�w���#dStj���h�&v�_�}Rk� �]W*����ۣ��/�rO�)�E��_�t��P�7����a��,�ݟ%����&Bn�~N7{6?��i9i��;�x�o�ϛy��)���9T���	�[9ۘ�n�Io �@��� v�hZu�_@ j�(�3�j�4O��u���ȥ-7'	���+�}���!���V)��5O�b�{��uV"��~d�3N ���r�z��ί�Q��#����В������X�nx��(e�s�7�%�?��P�IW&�6��;��қ_έ�E:3�=�8�꤬���2�/4_Y���ߧ�����׫D ��}ޠ�A�h+;��t�Ѳ�E�X@�m���	9�1nP�?�L
V=Z�����X����Y����W�u��x�x@Ơj�kft�j�	~y4���z�ex��.]t����(w���&��+Jl�����M�O��]R��q��R�ĭ��7�<���6pV%��������G^5Wf�M��)�ϬT��Y��2C�Da5Z�J@�dP=�z�33���z���2Kmt�m��k�s�B6=?b�����V�Ikc��&%V���3�H���+]��Z����%3���:%H�z�ǘ�{�A�G� Ys�#l#�2^�#ߧA棲���C[�N��j���� �NʃQ�
�����iO'`����T��{�����k�=�g�f��sfx-m*$�`�tn"��/Y��ZWE9�事�PGH�H�x���YP����w�n`Bt����L=�m�F���^��~�HHo'!%��49��($��P:sT�������L�d�͇�͑�݀���PG�̱����+���V����=9��t���+��`R_�R��zs���� �'0�`A)V�[�5��ZTd�Fi���������� ������X��^��|��e�OԱ4�������9tBy��f_j���T��{5��)yma���x���������s}��Y���f��Cp�9/ׅO�U$�������01ƹ�w]E/'Ӆ���ţ�H��U;)�4���b`�
�i���f��|�X�g��PX0X� ���JCم�tb��g�c�-̺g��n%ƌѬ���O���.��t��I����)!���>�k�{��7�h�0�ހjD^�C\��qx8�tA|�5��	���H����#1��F��iɍ_��YQ���A�L�^��`��B_G-e~����5���_�Q'��J(D�m���<��Yߕ̨pk�%����e���uoH��?���`�2���fφFN0�'�Nm:�8.@FP޾�H�wG�I�H��Lꋏ���}�y~�U]3R<66P���J��_���,�f8��J$��H��O��*�K��sL
��u�=���g�5�	���wc?�\s��h�K��4Eь3�"M9��������0�l�{��w�_ T^�t��LM�v<9���')�8C� �I����'e�f���'�|7����/'�WS� 5�P���YA������JU:�^�P:{�T1,�A͝ȒМ�(��$:�o��}��b�O�P|����`�I�<�b$��˕��qEE
��aM��77ш;�H4���)iR��p���S�qf��0��Y��+��W�F�%9�(C�ṫ_�t��ѿ����	��ōή��c�-QW��LR�x�c�ל��f�ƕV���9,V*p�'-��n2��݆�B]�	z	+�f�+�ޣ����b}*�	�=W��Z�=VSR։F��h�U�q��
���K�ߪ^��*(�?��E��{��ĵ9yj�K##"+�.J ~%)ZX(9��:"L��A4�$z6#C~_wwNBy`NK3G[��:p����Az�ii. ���V�͖2�-ZL�7-�R����Ou��}h��sYX�}���s�ˍM�����*�>t���Q'UP�a�\`m\�s��te�PJB@Bش$e�.'�i��t^d��c����\���!�D]w�VL��ޜ,�|���ׄ邗��{�O�h^6�+A
{y���\}]h86��U�h}hD�B�4b}�t`��8�MO�ֶU�������i����t)��R�%��Ғr�{K<K��྄��̦��7����jD�b=V3�9����l�p�2��vF�ЕV�k9wlT�*j���GA��p�ݭ�s
{���p�bX�D`�0K��Lu.�NV��C;�G�����Y�0.�ngM�'�s`|�T��f�V���kgBg�ӛ[�Qw߻�;nP,S:"4�p�6՟������	��<�t��> l���X��zx���ˏ?�˫��߬�$8D&|T��U]h+�R���l��]�>��x�5v~��O{s��|v*�Pws�j@�y,���*s��G�M|���snO�7Xh��ʾ����{�J������y�����[ <B����L���* �J�`.�Ǌ_J�.�����,�>��d��@#��G����Re����0p�@�1$$���h�^����a�U�.'�n�9T>�G�A�GSwi¡q�.���I��$/�? � ��i�����P�x>�S�$�z;�h�x+:_u	���x��������tb
�_�v�G�q�"�8k4P)	����HxUF�m����wO�X1Qb��Y������v���GS�M���ͼߧ���mJG�����i}-�"+|#9�����
�;+`Vn�~�>Z���l�WOn�.?.���u2�������Vɺ�J0�H�N�)"�����;Ds���f��9`�7N?�ЅZZ'�����n��[o� a?h�0�*������h�ޱ�B`�
ޗ�=��t�I���4�M�������k�ۉ-V�=�Dm�+qA��	��W��O�n���0p��K�/��4�������]��� �}_�@��*���1��5l*����Ƃ�&ٯ�f��.����*k_p�@,��ۉ����P�+�g]+,S��V��Q�>�Iqد @k��F�/E�'v�%�u�N�գ����9�c��O��cLf}��������ߞ��9�]���/�Ɠ�{�n�������~Y*������#ɢ�*`�D�㼔�����0��d-�M��Z7;�����ߕ�޼� �?��c��tn�#�>s����l�ވ����엞��Y�7Ȭ}5Ij���_j������D��ٔY����2�0c�޿�N��������|��]�ީX�T��RV-f�������o���#�ϰ�-þ��3�F�G�$�e5�T���?6�������6W\l*���*�C����/����|#��ߏ).{���>�տ췶�~��ҩ��N�ߊ8���3�5�g�e�8l���5a����N��i�Sn�=�ߗ��������+�~�0����=��3���ϰ�m�.����m�����ޙkn��G�r��~S�s�7R@e�^��(��ݭ�W�V��h۟��}��T3��g�E�珋)�8���s�"�mr�]Vd�|3ӇpBrs�)��q(���3o�w͗$9�M��F5=Mj���UG��8��������ًp����rox6��Z��a1�>I�r�I��,�Ň�����F����w�W-W���&��pO�zj���j�Ղ�$P��N�#�Adǒ8���AA��/� fST����g����^���<�ͭ��y����xT[5�S�TE�SϩVklQZsK͢���O����Yh�h�1A�UR51��HB�)��i{�{}}�}�+�p���k��Z���p�=�5�@�ը� u]Ǆ�LW&���t�8Г:�[K�M����$��mi:��ޅ]<��%6{�_��lȵÅ�f]r�	�F�qY	��'p� �.ߏ�~��}��ZC�;�ډ�ۉ�3>2A�n�����]#am���ƹ�O�z�|�.+�P�Jb.ީ��rH���Ύ���:7��Z9���o�o��_j{����	�_4B�gu����Φ>L	l^|��d�}��������>��@'�����p��yz�%'.���[��]���_�k�Y7�d�p��|s�I�XfR��L߷n�"��YꥶE�Ie7��n~9���5v|�e���:�Ӊ��9�7�K�/��O��<���/���#.k!��뻯h|��O�Pp�ܔ,p��喽,ʓ������� }U��s�^8�)����lqs~d��T�?�w~kOK�|�Y��T?�5-��d߼��������ѿ�\�%��
��.����(I!�g�T�W��^�h�e���������VZ�S�K�A�d���]��)X8^�2�,p��xWAA@�&�I*� �VzA5_�ۣϾ��"l�L6��T�oW^}Ex{l\;dg 6m�#�nO�s{��eZ~_�z}sƓ�A3�99��C��HF�S�u\��|�]r���﴿�h�$I����g�wc�m_�°f��-�eT����vR��>�_��ƈKm�oH�CS
�b�vssË}��3T��<�j�����[�@�Z|3�T\_�������f�� ���=9��Q�	�/�WB�D���́[)f�\�q�]�Y ��^�}�S�����)�Ņ�6(|���%��ϡ�߈+^ߦ�[������/��������%�V����@�ا�jt��>yr�V��$Ss�RUk����m��G3�Tm�ۇ�U�J�>����%DN"d͢?���KY��֟�s�FS�'59JSDX�<��C=�C����ӂYYZ+��И��	u�����E�A�o1�d��'="�������w����?Z������T���E��*�փ���K�Pw(��5'��]D�sq��k���"��]}iq�d��Q��k"��5��lB$G'��k��؞��F���fA���ڵ���OgT�?yr�l�=Ҧ����$NR"[��@ou����}����z3�z5�,�U���}���\�n����Jq��I@�tW��Ї��B���?�+Gy;z�7�+�Ԭ{m��cj��@wm���@������`���FbRO��Lμ=x#2+*�㇟���Y��&��Oٵ��͠~Zq�jt��уS��f��=~IS��A�/�=�}�H���hE����M�(�C�'������ٷL�� iZ�F!��[[��jo��e����j��Y飊dղ	W.)�?�������_�dYA�`�Sc�Uo(��m��qO�,�ig��3z�z��/V��m��TZZ�4?���9�U���$mhB\%wHD��%b��{<8�m�\բ'�w�tlpr)�3�����<�01q����~I�"���������%�v�τ��1Et���}W˺��?!s�����07�di3O��_��W���`j�f"ȃ���	�
�26�x���ʒ:z�;���4|�N}Ig"�=7��Y{^���+����_Ԉ�KU��9�X����.8����T�t��r�c���R%,�P)���@�5�Ώ
���m
��TM�uɹvpZ]�� ��⭍{Y�$��waV0`)	���ƒ�:X�Z�sC��s�hO��fF���u^}�=�6���R�I���¿ݤ��ǍU�������b�=9t�J=�v8HQ�B���O
��q�E���=�[ex���>�Ao��t1|��J�5G'l���]?���I���$u�����������������v�>x�@[���&[܂ֿ�9��mM����v�����9i�u�u薆�E=����~)���3�O3�!�hǱ{��䛥v6��z������%�%�����	�Ծ�t��n��E��>U���`W�p'�IuX�$a,U��)t�Č��Dg�����w�����=�P!K�U��$�M���F�Dy������>��=�S�I��k�c�S���p  ��#�oe��0a�	#L�������@�ܸ��hJ��/GН���c9 ��5@ôxH�<���8 �H����C�K�x���ֱK=]��'5+?^��џ���w����������DS��ScfD$�|��������;m�^n�aǋ�K4�?}�<�/���һa�3�Y�qs4w����⇒4�>���n�i�	A���zv����ծf�?����Y���W�x�6ɢbs��&7�B�V��A�oĀ�������Ɵ�Q��u����$ã��;�Uh�%��T�!
is(,@|��M'���ß�酐��"�D��� �7�y�\�3���J!�&w����Qu��í���Wy�v��'�!�y%����#�̴�X��c����>��p�����^}Y#D)�]����	?eR^&^ff���N�����6G��'�Oo��î9$�Y���ݹ��8��;\-���[%��ݳ6H}���a��Z\�18�^.��D3�lDP���Cr���ZkiE�sm�n������+}�䉹��1�~��0�����92������ <˾�&������ -D�7k%Z��L�#�E�����w�Xo��0�Ω�
=k�q��_1j8���D��+f�v{5��5ٯ�{\( �4��7�/\9����8�l������_����(�"#ü��EH�ϸ�<�V=<%PB)}D��,�$q��x�[Tm�)�%�mb��%S�Grm�%w}"W�v��ҙ*a��惘DB4w�CN�|����bSf�Q��b|�1�:m�X�|��n���יU��A*�w�*ujT�<S���ZZ#���=tu��*e�7C��hR0�Nx�4��&��e]y�x�.�f�Xӌ�<V~2f����3�O�Z,��-ֶ���L�6r�~1�m�m�}��s�暓0�w��M���ɾ��,�@*��b�2c�@[l�>Y�`��g�'B��rX�Ȣ���)�����/��3����c����/�kY�m�5�{"�-��>�Rf&�U	��GA���2�^��c��E.dw2uqL�B���T�E��hN�_3��V�k����[�e��ڣ;��Н��&�ٝ8���Z��l�ަj��JqFxt_~�ְ �����#o��&�c���v[f����s���1J�+�X��Œ>�SGrrl�~G�u;�Ʃ���D0����cE*���B=ټ�����!�C�X,g#�pawC���fs�v�/�m˄��0�� !ם֩V����\�;�a;��67�§�;һ�^G���'�a�,����t��n(�}��ճfN��#�,\��Er�VT
Yf���d)��O2�d�VM,c@��;T�Qe�f)ə8�2@�IJ����۔�*�N��8�;6�ؽ�'e���.	}�Tx#'��?�b�c�mx�|Al�����,�	}��"Zى�x\`���O�9���`C����������F�=��5��� )
������:����N��4��fcw�>�;6��39��Xw�J�����2�yy��H>�
�v�?�f0�W���������g���]�����f��3_P�1t�+ d���	�dk0ʁlf����"�V�L��~5�{�Q�ߘ�̼c��.�
#�D�_ˉ@j~��^l��j�����'�儢�5��^��$��-uc\�g�r�]����Y����M������P�u.��Z�����{���-�4n�֝e�ٙWtN��\��杢�9*�]�ӣЧ���ۮ�ƹׂ�w{,8{5�"efHh؇Ң2��0ـS��ݹ$�n�^��Z�N�H��
_j��l�XTk9��[{qKA��R�&OfN�[<WL�޲���r�+�O�1j�j��S���9l���S�m�����D��:�ݿSu��`~�&'��=ͅ,m�l�DC��FqOn%YS7�[V��p��x]��1���>�;�jԗ�;����Ѥ6�1��kUz1���qqCJNH%ǚ��\GK�	�������\�A��^�ugM 	M�����e9�˖�=XPM-�x���2��n>�������:b�H��5���2��՘��Y(�xԟ��:T 9D�*z�mt��+i�X��\uI�� z��ǵ8S�L@�'�btfek}"���ev>���XQ��ؙ�'�.$vDe����d��%��GJ
<%�A{Ĉ�I=��s�c��Ow�A�9��U&/0��CL>�,Y/$,�\���<3ݮ.�u�����?� [ u�&]װ;g��;�-��*�-sQ^�$���W�oHƬ�3�q�A��.�y�_�cD��S̘�U� �Ͳ�"LT��26���j`����\��TT�n�}���W��g��F3�d�W���pT��l{����I�OOhwM@D=K/0'���)�0J�4P�S�W!}�K�)Q!f��NBvO��<M�u|;�z|�nb�B��v��ޠ�m��{�D���y���߿��h,��?��Ν\�սy��Rh�t|������,U�������S08~�[�1�ԯ͐���?�e�x��.�̼_�'B��H���j�話��wm��4�WoG�v~"<�Wt�r4j�e��wU�Wq���ew�֗��-t� ���	��Ӂx��o�'L�j����<�J���yIN���{^��n�h���qK�"E#�I#n�(��N�Yq��ZGE���¢W_��n�y6��&QXO�q ���O�����*#uZ3�^T���wG����b趖ჱҐ�%��/#.Z����{x#��pb����kƧ����ݼ&f웋�Ђ��ϖE��|������3!��'����_Ϳ��L�;C�Ԍ�1�=z��t��>��Q�eN��͢����g�*Zգ��1L�ϸ:'\o��/,��ll��b��DN\i�0Ox8��	�H�[[�3!=% ��#ѫ��^�-(�Fߜ�Cki�B�o��I�E����u��x�E62VN��%r��Au���u�;����L���2�3L�����r��TV$!�Ϻc����0O������{رp��v�ʭ/��M\�
���;�V��O$�Tm$��Y8af��t��h�'<"(�M B�M43u��d�`�Ma��R��j��w�<�u��G�=(I��셵?K_n@�v�;ʉ�W�D�j�|b�ݖ���.
j�:�A�S{�����N�o��q�q��*`��h����RJJ.A�u]�hB����z�f.d�s��ctl����z�3l��a����Փ���eO�'��d�@�Z��3
PT*A����f���e��:\z�$�DEAQ��WM�>�O<��Cfm�wU
Z����5��Jm~<3O�bt���$�N�o��6n��6��0��k'V⶯H�*��9XW�2��g�y��+&@�F�%�0�i�e-��R�]o�?��&вB�e`(M�m[*�w�p�涎=Nlfp���dt�.ݶ*��p���ԉ�ӆ�@:����4$��tL��R��!�q�,x���d��ڌ|�d:��`�5y29����5qq�5��!�Yd�7{�v	b+�K�|�v�c����FTZ�m�#a�4�/_�e� �/#�v����a�P�ѕ&t��l���J�K��!j���~���k�������5w����<�8��`��� �	!vyA��,�d�.�N�~=J~NS������dr��H̺b㥟��p�?��Z�|��{Qݕp�bRmbo�+����~��+�B�����M=��Q�.w��8�T�y��_b=�ۋTer;� yC��h!(V��f��qW�'��[K(R�"Y/g�8o!s�'5��Ѵ�(9<D�1ƞ�%��,g�Ɛ�F��~ff�K�z5�����S+��>�~J~��x�3���T���R<�Ee��G
5�n}
bo�.���nFq3
��[����<�c���&���a<(ry7Ztx��y���u�nl��-ѷͿ��
[���ʟ����-��4���̱%�T�*��%�f�y�(�$�/�a�u�]������Pza�#���~m���{�}vV�#��\�_x�:f)��f�L=�0e��nKD����|0�js:ٌ4p6C��ֆ�R-��^��Z�fyGQ���J���jf�F�kQxC�Aʓ�/�8F9Ue{l?��N�����`��_���;WM4D?+ׅ	d�,��2�=[�fr���� �U���~;ZE��%���)4?��V9��)��.1+w��8B�WHk���=��T��Ly
>Ez�N�r�F5�W�������H̥8�"L+�Y:z�Cjnxv��ȷ��1En̒K��r�+����2Y���ȫ��ayM��a�mwXޚM{�-�`b�`�c���2Эz?� �"���I/j�_�L+�u��f\�^�T�Y��������0�|W1$B�=�HA��6��TB��J"�١Ö@KI��	x�L���Ή������"��A��'t�W��2*v���IS�����K�߁A�]�b	\F���Q1��q���e{��8���:�'���c�x�g�� OZK�$�Pc�r3��2j�M�%Q�Nt�Ԑ���VO�^�j�Y!Vr�(@�7�5�����[f*���
�����������m��#�u)�̷-*��R\,� �-/a��h!6�jR.%�9��q�³gVC�b��[�za�]^=V��|��a���D7�~#)�v�>g.W��cl.��x�lCﲣ��k�<�1�J����i�G����/�{8�E�>�S�l\G�y�p�G�6�S��?:�����O��C?49��}��1�~�f$�AZ�c�{3U�r�iu|k��qc�(%=�5����v���S@�l�'��PK-Zk�#˳��fc�n��+�)�FN�I��:��3W�n�z����E��_�'Z�z	e���i^﫡L�N?��M��P3H�VRUM�؍�%Ǳe�r��+H�k�N��˰��#FO1���-�?���jo���}��:_�S�^���:xC�_Oج:�]�ٓ��g��r��,�N��^\ꞥDН��a����>�D�N�/Y��mG(�t���nnf_̧���堈6�娲�����F�U�ҞODVI	"=����W��NO7�t���;M&����l� �󁠤w���C*E�{8n�]��Gd��ΡWA]�zT���a����+6MCm5�8k.�W�?��_�~+���*���ǆw��J�������\'?�":�fz՚�pv�*5���#�FZ	�.a��4	��gR��v3	+���t�}\�st$U0�>nWC��NR��ݶ��(��Y`3H��&�Q~��P�q��C�]+<6� j���3�#�Ez�'����#����~>�=ȃ]�ż]lB΃@f���<0��ք����K�C�W�<+�_v�b�ؠ(e� �Vt�0�_"]"�߅}-�[�[l��zڱR��IG�m���H�Mqï���Ս�I=���K�W�1�fF2R���-E�p�g�Q���xP�ɘ����Vɇ1���3�on�s�������g{�p:������pe�`#]�p�������DT]��)2���L��WQnE���w�Hc.
֕� J
�ftn�º+|6���� e^��qX�9lq6����F.�Ojh>�I�KU[��u�h���ӭ��ۄ�g��q�Q����Λ-= m@�eη�\j��w#�C��nTx��>��T!��Pԛ�Y6��_RD����^�bH�p_�7�1�O���(��q������_�H������\Ō�Fz`~+z�Y�֔�ȣ���-@���*��]q~���<����߭4j�m�w�Q���V��pr�S���߃�� ��<�i�Y3k�='L�X$d�{o�Dy�݈5���cI dmȷq�2J��"_&�P��@1.T���[f�ܵ�������a�G/�M�BZ�C�q/�r��,��[�qyǂf�*77;��{�`�tH.��`ڧŃϓ���_�8�P�zY�B'�6J��5��M�J�A�^Oʋ������(�G���J�Nt����k��U��V�����(w6�Պ�z�w5SQ��h�I�hV��1�p�d~7;�<�_�du7�+ �,������uI�?�z����������Yt�c"l"'WS�ϝ8H5늘�	���HN6x���dV������-�{� {�pv6%����8kt�p7� e5�W��?��z�
�������v�������P��2�2[�TA92��r!�p8ć
G>���#=��_������OZ��}��~)l?;��|y����a���u����(�q��K�ȵ/��,A� ߙve�'@E�{dۿ��4��&4��SSM���ZZ^�w!%WL�;������؝" u�$�H9����햘;�
�!4�eȚ�3S!?�<t�ti8IF����`]:�>	�3��ǖ7l�f�t\��4��~��N����w�r��c����_�x#u�_����ɳZ��I��b��ꄖ���vba%�Xk�����tu�J	�-�h�٬ow�7j���o�qCah����)�H�<�]�Ш~oCU�z�9�o�$TQ���C�;�\�(L��%�ǖ񏤽�i7� _~�_��y�R�cW(�b4�x�;<��� �:�����=��Tk�>� ��/�F�wh��[��6�81��+�5X�H�h�u�I�Ѻ�So����Yg����V��!VkK��)��~��� ?�ƣ~�� :���%��>%-�+�P�-a���0��	��G���J��_�SG��l����'0~�R]�(u@m��9{��EN<���������؝���ME������Y�Cm�_HB���"V�I)����_,����<�lR`c�P�~KW���H�*$*�f��_� �+�{NqWJb���xf*�����y6~�)��i��`AЅ���\y�"zQ�# \#�,I��Wچ�Ӯ�����&�Rq�˼K�oU��Z����:oFZ��\�@�|-�k�b�`��MtFE��Y�K���Oriƿ�o;�G	NN5�y|*Y��/�p���7EF�	�Ǟ�=�$~�lYBm�_�\G2
�p�<�mnϮ,����St|6�s*@k�����{�Wbw��[F�Z7\�L�*�^PNg��.���F�� �E�:�e��A���2z�D�di� ��a���rlde�:�J#��h���"Zcy���P*�4Bi@f�����J?���Ķ�bBCw4�G��/���f�6ڧ���$/�N�J���Y$K�Ѥ1�_��O�U��;ן�k�e�����iD�|E��J�BJ���*�����[�T����>u�ii�0xmR��A=܁��<����s?4�TA��D����c�X�Q[xr�VUl�h��"��]?k�kM�aC
�}(�V�J=̚(^]�/$�R����C�6�Ԛ/Q��i��Y��{Є�!���ΊC1:9H�>�����!l���n����Q�<\:���)����*�U�+�����������6&ix��9(����qC+L�΍�Uc@8s%�T2v0�7�A˩���̹����`��*V��Л+��VT����^���0��.٘��,0�P�4F��q�ИF���O��S\�/ږ��L8�V�Q�9�/� .���rnqo��
T��e1	"��Y��_<�n#�[k]�>.��>vV�'���O� ��&���-j�|�Ρ��5� �@�Re!�z��+`�*[7� (�ӄ�Uۏ����JrۆL�@�oR�}��P���#�_��Qб|�X @�>�;$uW�¶\�&uw�0�q��9��\]N�K�⎸�A����87����� �X� ����z�t��zS�D�k�F��_�PNe
i�g�e^{]�Aʽ��0,:�|�ʌ���3�h_v��]�ê���6Sd�)�̵.�P�y���sIy�\�1�x����A`�a���!���>'��4r
bЖ��>S-�}��H#��ز�z^�?^\���q����C����o�}m��ʃ�џ�.��W�[[��,Z ����V�p�+������Қϗ�Z]W�=�,��_��:>�v��0c��q�SL,��G�q��5�YdE�O�����|F�D7n~�P�5�W5R���=�9 ��G��+Ud�LT�? �{xp�q����HQ�m���{-�`���s/���SJ�}E����g����>���,�7Ԥץr��#4�-�����|�j���sL���GO��f����󸨭f��f����ك��ґ�JM���vs���ʜ4�Cf5��Kп�"�)���@��i�*��(;"[�(�S*��L7�ۋ��.����e���@��e�y�� �^��hU`"�1�����	&�&ڣ����/�Fq��M�)�׺��ҥ�ʉ�;����om}ǆ�e̓���j�ϴ�G�����2���x��k��L�-���T6� �����<O-�|lYr�+�'��9�]�R� `���Bf�*��!ߣ?��
�wy��{&&d���\���o�Yp���bFֵ4�)����zs9�a��Ȋ {�c@�{m�~4�,�{!�ρ�g��x��A�8���ep����'swyr�&E����-�@�[J��B�^�V5p����5	���UB��G�!7\�]��5ֳ�|�@�GY�J9�y@�K�1^<I~�y��36qSS���%Wb3� �� "�1Dn�����ח��J��D�w���^'�N!ڢg�K�k�&7e��o�풫��9���)�R! ���{�E�yQ���Si�='6��i[tͼ��H��K@��K�m?rEma��}'��,/G@�࿖�p��N{�<���i�SX+({I]��3�s�H��e��G�/f�W���H���xN��y�G�^D��Pv�z��$}#������h"����j���c �8:����k���Z��|�]@=��K����%�����`��N�/~(O�Qt�3�R�Yo[\ʲ�![�B��:��d�83�Y�4��T���LZ�et���@����� 2��kw�oq�0,J���g	�0��u0�0���^�i�˂�*,����+���H��4	��ACz�v��X�ir�?�?��ȓ�F`|H�g��?�{q�{��G�b��;E7�^m���:����G�
�4�/(ؑwN�f�^�f�w��cU����y�ds��G7���ݏtԞ�N���WSi�p�z�r'��J���t�+?7��M{�#��h�ս��s��`���=r���z-H+Q�2b�~p�*��{�����L�?w��.q��.g1�A
���p��*['�]ȓ>`}�.&��7
��@2��4���8����쯐���#����M��z{qhI��Q��lL��"B3����t��:�ʝ�G�
Ƈ�-���LF��kDq���lD`SiA��f���~��������;��}�лY��zj���^�%:��F����z6fBV�ٜ��t%�W�[����	� ������J�!b�/���������6m!���N�=� �� �{^&�v��� d��QP���%�	Ɠ��%o�ςS
��؝�����������JK�edyY�GZ�j�XiS'v�̣p<��=����>�tA�'��a��E@�~ځy��4���>a)���b��+vB���p��3�T�W��E��Wm��:6p�n�+�t1'Ux����"�����&#��9���v�ٕ?3���N<)� 6j�)��?�-�o�
��|��N[�G�����!��4�D'OS�"�t1�{�D�S��Ʃ�B](�xf�г�X����H�q���\/��m��D|#╉ޖ����N6��`�!�.>�/c�S4+D���RXA���;ςYd�7��X�a��_;�=�h�3�[)a���_%F;k�fL5���j���;�~i1_������<�=��#����gv����/$�@q���κN��@f�63_g��L�@��|����C�.��IX�n7��蔢��j�t�h��`<�!����������՜�;�.��x�2
�0��\h�c*�zw�h���p��\b)�~q��4�z����VW�^���ȅ��'m�MF�{�hi^��b?J��ڝ�u@�w��3�}}0��	3�T�m�g�ڨ�֞8�p�3z;�����xS8Y��2�w��0�a�oN����p�Ei�����Y����ɨ�1�e`��m�>"ec���}52��_�\�z�Pu(/�Uک=Q�o��]$H�Gw�s}�x9��<�I�j�w6��犢�Gp�3T����.��㹘���EZ4]gY�� :d2�{��j�n�~������޵v�;��@����.�ğ�S8d+/I"�Q	R�C�!��w���H���CX���f�^��ۏ��+�vI�3�ND+��t�kj�N\3Y�K�����v��0�/i�4����AK���8H-�d��@���Y�e�g�]m�m9��б��D�?S�M�<�
u�~�a��H���<�R
5׾��i�C�褵R�*��F�n��3e������r��Dۗ�R�ʐY�*�}>�)}jL��S��Y���Ԡ�@w���u��'�-OR͛2�H��@n����(f�d�L fƫ�5C,qN��5�ng<�W�*1 ��L٬�'/��-�ႇ6`���j���������Z�&�!~�~H�C/��x���w˞e͈{����/%�>͠�OzY!���R#CЎ.2�{�5b���J�9�X�ny�b��.�eu1��M��~-e4<j7W	e�i�[oK"T���P@��ý�X�r!��nM�h9�����KY��?��L�f�CKߛ�z;��������[ߦ�J���Fr���.�z�	����m=�#��v���Ȍ�m����k���y1����9u��V ���zr�-�G�tג�X�Vʍ�0�A����]��^�
)�?�蕧[�_hVwH/���
..4,��ڳ�A��{iz!۩�Gz�![Ť��c����{k�`a�M�hZy�t�<nu(d�UC�����p}�g�ُݵ�'�ζ���z���9v́w_��R3�]�$�Pj��3�������пR��{@Rz0��E�����xb�ӎ��y:S��j��% -[_Թ�ޗ�UBu1�y�t$�ݷ���� ��z<<5v(ǛN�f�ڔ����O���z�Z���P��uO��M˃�L��ol\	S��z��f�����[N2ʫ�����J�R�U��y������- <S��/�a�153qH=��v{�ͶBݦ��j-��	 ��b�&#EX�R���T����'�O�*�y
�W��g�	�y�\X[�|�(ң~FIUYF�9"M%s6%���KT��W�*�
`��-
�%��lci�X�܌���:��C1]|z�����J�$`��W�]8S�vkx��Z�s���u��$Y�(`+I�!�����T��1C��f�"Q�Fu^�6�Y.��y3�1� ����Ol����HZA֫(�D	�d�L�%��p�f���$�\�]��[V�W ��+6�&&4��+@1~�Z��z-O{>@p�s��VK�v����y@�_��zַ���6B&��TV��焔��Ho{�G��%JU`Uٰ� �̙^n�(�-�s��/]�J)����=�Oq}��A��7�<3�8��rO�HaPް��&�H #zM�Ғ�%1����c�e�=ڋr���x �^�a�w�ә��j�`3�N��PK����0�{K�E����"�(�F|��t	��λ������,�H����"�&KeI�%��`�Ab'�xdL=Su�V�G	4B����:i����GIU0��-�W'Ҵ�SQ&��
hֽNhF�J�@�;��ktR��k$�����Z�0~n���36����sB���Һ&Cz��t�i_U�h�\Ph���A�C`�<�V�Ԇ��{�l�qM21�~n�Dn"h 7���6x�i�NШ����a�$3?����H\�	Q���$=Q Y�A'%��h��u�h���{7K�8Ԓ� ��T\��S3���r����� �gÊ ���U:�����}�i�$�Bl��{���ֽ2z�
vA(�6��/w����E5v#�չ#E�����Hu�K�H�"_ix���[_6�nN1���6PU;e$1�z0!��x�9��$��b��}�/�m�n��/�M�<
��Q���B��ϝ�}X���i�\r�^���V?�7pJ��5x&���F?��ʘk����W�j�/��߉lH�a_L 2a����>m��*1�jN�m~��z5���;��0o����ԍ�o
[��;�*��#�Y��a�o�"/�����oQ_�i"�x:GRGf��V�����4���ɒh��zc�A㺎�����ڣ��f�ߎv�y���~Ot��]�:(YE�D�9�AZ����ᾡ�?������q+01SRd�L���}�N j��ro2��^�G�qX����]�z�1czŻ�Ti��Zr��F���vF8~�/�5F�cJXF�E�1`��4F��<�{�06 �e��E�O�&��o�ɢ`��ř(|�GV=�@���+������P�)
ڹTtL�X��^+IU�裷�ĥ� -Q�m%^�����P3���~	QO0G�h��~��N��9u>9����e*sc��f�H��[\LZ1�$*Ze){k���&��W��8㤚"y� �0��h�)�H:�cV�DP���4�.���w��x;�=��]����=x;��RA�?�i���;8�!fp�������'M
4F�/.�i{�+�����T/�I�� ���7��Ց]���kc�w�;���?i�\M�5�W՞������q�����f�=�X��nV+j�1�F+�d�B��Jco����9�����v�vx���2��� Q�`��=V���ܻ�5�G[9���b�ƀ����p��9��a@ּ( =���v�e/��l��6rZ��4%��J�3JK��V�A�Am�RV��S�ɇ�˜���a��g[���_]�6�f^��|�b�a:���v/�`=�c&J.��9SC}����(q/�6�ꠜ�R����a.D]C܄d���c��I�8R9�P���Pl/������C���@��.��[���H6�$ݲ2������%H_0,�Ŏ��GɉxY"�w
��9�@�s�j�k�C����̘����>z*ūξ,��y��j�G�ι1���]}[ߺp����s3�v��t���^���������w�ؖ���NN��'(|^��<p˃�f��F)�т�+l���)r�
c�����6���Ț���[+�y�J�m�\i�����]Wf�M�ׂ��vJ�(%V��{�Vrs�M� ��v��dm�m�0*+w¨���ˤ�����8H�����Ҟ~f��7Y�Ǐk�����^��-Rފ��%�VhJ�v�{�{\N+K��1��_Jv����p� ���Q�c[�toA#z�b{d$�wi�>�Y����z�.�G�3:zil���O��X+�&�Rtu����Py5��E��F���4���ww��}��K�X�z�щ��O~��d�R�rY5)�>�A_W�����R�Y��<�a�E��:Y��zsuh�şl,q�`I����T���b�7�ʖ�=���A��n+� �h{����>B�푄�y����*r�_�
��Es�F���^����y��ɺ7-��>[�Q���Յ�]&�f����6�ѽ��̄�Pf¨������S��d.���,i�j����f$��A�<�6'v�*�㇢v��D�F���)aV$C��&���QqV+���_R�:j.hyN)h9C�=��W|�����Q�U�	���W@�璞ROe�J���X�����+{���ґ��_p���\�1�̝�W9�
+Ujp�.�����9�1��;ڵ�ԁKu���y�o93�Y7��:ܘ�<W}�Ē(+��n�Å�wIl���OE�Vi�^�b|������ܜ�Įy��΍N���A�_Tk�*����bV�R��Ƒ&H�bɗ1屒�1ԉ�#��d�i�W����xmף�(��I�]ܖ6t�s%���T[�h�U�����[|�����ֶ���c����ɛ��~A��hVt�\�er3hl%�LK@��e'��;�P%���C5�@��p�x��'��;�]7*����X�$u�����/3��˦��~�t���y�m(��l��d�H%�M1�k"#�+�o��f1c�Ƒ\�1L�|.��Ws��]j'�K��"�u��{<30�8_���;��z�ݮ����q�"8���QT�K�>�)S�a랆�̾�~ZM�0lTi�AC3�$���\�Q�seWK�L+���ԙ�e�Ɏ��96}�!�ڐ?�F��{$���~��@�(Q{��z>�ꮊ��f���?d���x(�\����F��fdg�)��9�RF�z�mv��5�d��c+��1%x	�}����2������^�S<��?=/-��K_Mk����Ύ���M�z���V`|zBZbxse��ٗW��^ҷ&T���HĉW
[��[,xTG��0�:��!_]�Ç��WDU�UN��@Ȋ�P��>���z!��z�b[�l��� "����v~^��z���0	�ʤ���ƺ�ݻܺ��Uߡ`cc�\n���/�Nr�z�o%Œp�h�Ou<��w��w�>씽R�͗�r�lw�D~�HT�
�!F=>q������N/5&����+��`1�Ȋ���V�Ni9(է���2L�v�f{���;�����q���
RGP�bA�"(]Z("�CB�0"HS� �I�t��PBI��@����n��������keɊ����g�}�{��t��d�j枣�i�V����&��O�\���+��+D�C��,��^ee/�Ra ��>D�I)ڌ����D��/R�lqr6�\����[����&ꚶ�Z�a��V�� ��و{%=�b��Z�'Gz#ON\�s+c���UyC��w7#e����baE����P�N��_�ߡ|3l��E��:NBmH�7���:���/�?z�{<J��k=�yw]܍9y�P�,J�5���?P�'��3 �i^��{��Si���9{X�@S+�4k��t�Fڑ�/������lEQ��������cIeQZ���*�\��Q�v\�x��
q�^!���;j�yz<8o�"��N>S(��r�|E�m�C�����J�X1�����e� �ܥ�4G_�w7s۩kG�F%H)pW�j�ޮ����&��>�x��J(�li�?��?Í�)����!��L[o.r�yG�����.�&������I������5���K��y�|��?a�.����몘q1J`��M�J�n>Ӳ�Q��B�Qm���G���d/�Q�(�!1i�O�X⢒/�s��VQ��E��K�(����/��X$��g���]}x��V�og�kF/���]>�P��u]n��W��P�� ��f���qn?u�>�.j�ʹ��(3�8)I����'��� @���XD/5[f�e���W+Jt�cJL.��W������䣸��O�xY��ᦥ��a.�y��P��Z���\k��J�>[���!{y�r��EU���s�u�~���u?[T��,
�Q�*��ل��h�����9�nϚJqf`��P0��>�!��@���9C�>H9�`V����)��4V4猤w�uF�Ĭ��<X��D]�U��vs<���7�GA��*�}r�C'�����c�%�4��C5��ӱ�=�se��.j�I�e�PS��!z�RF�t���,Hg�i96�W������i�$�Ѷ���:^����XdGh��=v��"���w��t�K�ш2��T�)1
Y��F���{�ܼ��H��3��
�Q�1��}���`�k�u�|��4B���"�K����L�N���<�ȁZn��f�pD�;U��õ�-�!:��Vݗh��?pr�ߟ�Y\�$*���w>P*���NQ�1�_��1�q촁�)DD�p�6��<=^o�`�:���@���ݿ-����`|Z�fG���s:�4��� �i+q�,��S��V�!}Z�����}h�i4�x�&�l��K`�^�5.tH��ѡ��}���k_tb^���;�y��ie��8NL:�wL6(��֍��ҀTs��R<F��.#iN����X���q8+���������w��i��?��*�[�}PR��q��g�������
���̃zs�'��Z4�z�w�_�@H!je���A	e�J�탇��ɻ��G�L����S�1��Z���$'3f���L	-��9��c#�����n��.z4f�q�G��6�����"c?5đ7�5��Ke�;ṉ����u��U�Z5�H��27�9���,�����J��@������J����×y�xL�����]���vr,�.{cR��渂��ī �^�tP6�	��KY��὇�	`f�h�(�f�[s��M]�yFy�f�V��"z�$ZS�^e2Ҏ�����2>y�0�Z�ir�x�n|�]�}��#���sg3��둲�Ϊ�!K�����MZ�)�1f�[R{is�IPCPw6���J����f���!���<I�ؙ��GƇg�? p�q>��_kt�\<��]L��q�~s}B��KİF�ȱ��������F=���K)�ŏ�l����p����u��vW����R�?���3fGn�i��S��G���ڵ����|� S�*�P��A��U�~��D�l-"�d��� 
S�X��~�_���pN�������2J_��;Q4H�u�W�/��}�<�kP��N���kd�Ol�Q�m�\X�.�b�x�����͵7Fܗ��)����,dʹ����X9�%ݗ$�c���v����Y�����`�wJDw��;*���S��3'��
���d��Eg����߄g�|�b6侣�!���'W���8��A&]���##�4k��ٟ��6.Au��H����l[���+�<�@�Q����^��F(Ezb��^��d3�X
D��7i�!�7�+M��'��/y��B)>�z�<1j,��p�A5�p�I)���勿�����[u�u��BϏ׸�\� �Zף�����8ZWv&�'�g_w=3�?�����B�tu+@ �����2��U�ox3S=���d �4��0��=�2m͐Z�V���嵲)�1��t��.>����ס�Q�܍��������N�,�⏦n�S%��(Z�����Vv/za3�����q~2�I��J{�9"8�`I�0z�[r�}e*��R�f��'�'/a�o~�i��z\�\��tM꽪�\s�x�h�� ����2Pk�K+�K1�ܞЬ)�Va�Prk�k�]#��	��Y�)i�$�jJ������`�i��J�c�^"�8����זi]��I�la�T~w���н/`�W�f����U�^��� �7�׽/� &7��I���i�^V���k�U��m�j��!6i����71�?�5�Ѿ�W,��i��8��Nm�ں�w9;ưA����������[ d>{�c�5��8�m0�A��Kz�'�����tլ/sqG�J}�n���@��m�ɣ�C��ۇ��؛�_u�Wd|.]z��=$Ӕ-��q�r�%Π� �z�8ݒF�[��I��uh���V��	�q(+��;e�hȈ�:d�:��wI3��g	ʷ_u�[)C��a�"�v�s,G? !_���z���9�^�zUL���.����O^�0`�l��ܞ� \�BX:��̬�ѠO�h�ͲI��eR��p�5R�DU�	�d���:��#SNC�����,q�*?f:\c���n��w����_<�Zd���] �Ru�@�ߺ�ӵ�������r�>13��Ǯ@����p���њ���N�'��b����z���'�����i�JP.��̨����5;��H�I}P�����{�Jځ���t-�ı��3tM���]�;���F
r��ݍ �.ǘ�uՉ�D�"��s�c^3kO��6���a:�n�>(�9�JR�t���N�Q%U��Co�h*����n�Lrܨ���@�K��3�X����ҫ��<�;���}�%�S�$�������]!�/���}D�b�j�e�+�Q]Om4ǟl�O��0�?b�����س�49�\�l�ޒ�?\]���:��������ջ��^oVn4+`�B����ȷ��z�Xc��_�K
�K��^����f�j�X,ME`��%��	�:�)q����4mᵧ��G�����W~�՛���"\jZ�����o,9��*��`S߆
�Mf"F��O�b������zL��ͨ�*���/��]���Wb��}�W%V���, �ߕX9�) ���A9�K�N5�ĵ�O�a�ٌC�51,�Z���1%JZb;F-��S��	�˼�� GF�\��g9�|����ËΜY:�y=L/�6�{?�\��=~�������<ﭜvñ���
ïUU��~u��*�NT���ri;������/b������P���ZV� � �[�O��>jN;�P�Ȕ2�����(#/�o�$q`{3|o�#26 >��ma�	N%���Y�(䫋�ah@�c�+V�\�gb�����o�_��j��?~T��	����?�/�6�6�]�o���9���@yo�oh��CQ�G�@lt8��ȑ���A���ʹ�Ъ��X�`:��9�}W(+�Q��$�>������ͱ!�:�6`<���e���_i��s�?ڀ}�@�|�$�?jF��V䮑����,����S)���r�?��Jw'��U�U����Q���8W�N��&�X�G�ư��m��C}*#�K8�ssV����jUf���fc�a�-!�Ce�;DGJ"Y'vW���.�rhX�������^���?��A	�{A�厾T�
�O�����u��όK.%��<)!��yZG,b�h��у�����f!\hZҖ+ХV��(�h�w�"c�M_�aw}�CUT	�2���F_Z�.��ӌƽ�yČCE��R�w�"�_vm��'��g>��E�/�}�o<��Y�A�!����Z�/?��hf�`�:�<���| ���Ŕ<�iоC_S����OT0 9[�����Ip�\��*˹a@��� \@k(�{|:�:	ޢ� ��۰��{�=��dasQO�~	����p��0+��P�22��5�7@��g���{������O� �^�Zyp��0��L���?�,#��*?� e�S�,sW"[�,9Rf{�=d]����u'��fݿQz��l������p){>e�X˥6o�E',i�6��(XL-�W#�x���zŔ�P}�]�6(�޳}�n���W4o2��\��ֺH��WRc��m��$ ���Q
MK2�%|\8eտQ�}�)Q1���zԵ�2�>�8��j��z��^1}�����2�eʹ�7�.�qڟ��M���dյm��� u�)�����a�M�������=����_7�b+JWh�:���r�W�uP���7U�w����� CUV�� WTu�愈w����	���ܟ�N^t��c����s_�P{1I��~�_���<)i��6�7ȧ�{��h)�x�U/5���?�������1w�����n�߭������������֓l�O�C�K�Y�:�!
ލ3�zqzEg1^	�������x/ �v���x��g��f���N�{+3M��vj��d��o3ٲ1�W8��ǆ�$+[O\�/G���2NW��\UK>ET��C7���?2?��0,l���Ľ�8�w�(*Ų��vW��5�W��M�/�¢~�ňdۧ��D�o��$�G[&=̔��h!�-1o;ۗ����aˮ��&�k��Qs{�V�`�O��p��Ɵ������;��#�9����t�����W@�/��owH~�p�x��5��%v%�3zg���A�6Q�SZ&t�����qWY�[9��W��Ų���B.ގ==n�������)L:&��Q�����h�z»�h;Qּ�����;W�a��m�QD�T������S,֦f�����%(ne�*?��a��D�\�my@2Y��\#�,�lu�������jWŐM��#����H�����D~wy�A�$���FW�_�(j�`ߝ���@ݐez���Z�kx�\ڌ�8�Q��h�\��E���7���92�6:��)����������9E���P���Ĥ��\�geAtX����i�������ZnƠr���`���g_KI�3�t�3�ҁ��]dr��ޠ���y��]��H,9oL|Y���|��|�e9��"'1Dw;�;�8��G(%W���=��v��i�*c;P�h�I�\`y�ܬ��s�gl۞"���ִ��HO��~��ޜ���YU����Z1c�g�瘲�����D$��]�Z�b
�b�~��t�Q�d�B���f(��HC��xGQ���	���F���\�@?76_^��?��>N�q�Kg��m,Ҷ� �<"�R}������o����gP��F�R�ҡ�����꣭m���R�Wá���\���0ky�H��V��e Lw�ri9�)��c�3 �-�����)��W&.J/�s�g<�����Ыls��<�1\j2U�� ��ņ�7�����N�N����QwHoC?��zC4o]�:�zk�=�<zGٙ�q�zo�}��Ϸ*^~������KtGb�&����v�Edh�%N^5��U�k4��M�Z����������f���)Bm�	��O֙"}U%�b�2��k�ş���Q��h��lu�+=5�c*��@�T�'�2C}��J���B���9F�AHZ��̈́�_�=��{�P���m-g������EHL/����5�Ǻv b3 ��Ss�vg��|� ��k|ʛ��N��W��a>�J���c����p҅��VS,ϵtEx鞻2��V�_M�{����}���9h:��ל��m�%{�WЇ�
$��:��K��8�@�#>6Zn�w���z2��'�܍�5��3ф�EE�[�nI��6{J�7�_o�<��-����T��j�����jr~uy�;�૒*�$I:�O���E��}�TI`�_/{HS��p���2�������K?����I�����a�?N���;	�7�����������@G-b z%��D��G�p�Kwg��$D&��_ ���7s �@	.�C7��[w�/wQT���w �FA�Yo^WۏY�r�d�C���U���S}o<A�uD��ZB���g����!T9`I�IR Dz�|>�����[�h�*2[���ϙ���*�o��e34�YQ�)�.", �Xx6�*8���쪚"��K7= �<M�����%6�E��y(x���rկ��Ϩ��J*ו��t	|kJ�P��2��֒ɪ�QTdÜ_�ͪ�X��=�1j�2cC���QXS�����?@X�qEOI��j0�|Y�W��Ԍ�q�Q�S���:f.���Η�'v�[늬4��Us9(Hp���%uЯ�-�\��s	�S8e#>�	t�_}Gn-�gQ����M�b�|Pw��b�@�����n���T���#��d��J9PG4����e����0�G?P��j�X�'�Ĉ��x�i�}��(+{����3�xi�-g;�^�`<��q��P�?�F�V]�,�^&ל�œ����\
�FJ��MO�ߔ�u�u���z�?���ܷ?]�AYxv*��l�u�S�x���2W��E��r/[�d &������Uwj1k��@�:r��#��$�������¶䭭ETz���̓���k ���gi_��~�U1[�Y��J&$��Xi]U#6��
��͆xw2�Z�^��)r��"�N�=�Պl�����X����嬩�t�H���V2�,�޽��f38�Z�0�R{hX�7&?��;�����lFD�W��J :���b6m��4��R�a#��=ee����ѧ�.�h����I�C�} ]M&�p~���74�G\7��|5��n�� B\j�PSESp�>�A_�_� ��R���pֽ��ՐGa���W���$$��2"K��n��.�����K��'9���APa���9w�2&�d��-����Ɖ˧zoh�$R�����&V�pKbR�E��l~<F|�� ���N5���UHH{#��#`���q���XOm�:�V����Z��not�Q�Q�̀���!�ŲKq�����j�T�0�E���Wr��*!o�z��/;}� 1{���u��#:��s�L$tO�֨aN��?����=������Q	�[˛�&�����n��u�'�I�m=�)�Y�K���3#&F�댈X��Ӎ\�-��^��uC�̙�:iRz��8�%p��30��ev�~2��G�J{g���y��_�s\6I�t�s���_0?��ڤ�F!#��r��Q��Ɠ^��#��sk��(�����}u�� �-Ǡk�5�tE�pB��7Yf/'o6dvH2�����i�]M�uJ��P�)���`:-�nꭽZ��wT����URo���MT���g��f�=Z�.1�|~~���nq�b��Y��g��
���'2s�s�r�o���&��䜹�#@8h��ܺ�Y!��J���K���3���`*V7��}^�o;'�5�RY����N���Х�:o�Nѵ��e[�����R,R����w]?4k�q���O����_��\;��"q��5�߇�z�}qJ�Ѐm3��t	/c�Ύ��hG*e�g{�T��2A��7��')E�l����F��ҴkY��4����T?l
�q���^��#���6�t��Kw���s���ً)	\��J���ye������A����(H������d@벇㞿y���9|g�y�!V�z\;}s��"Z�'�_�|���_�d��S�,�	���&M����y�D]���W�/��M&N�#�fZZ���R��Ͻ����SJ0��m��}|�_���$�6�*�W��rC-�$v�r��A��Eq�>Cp�`�����K�T
Rn��~�a�3�=H7����O(Ÿ���rk�f2||<�T���� ��!z��a� �3�_�$8�s��$i�tӧ�D�hx� �u�A?�'���a�ㅃ��W����f�%ۋJӞB"��^�3��M��:��\|�U!�F	Y��)h?�l��3�3���%M.s�Ik	����0��8��U]�^`&aZ*�{�cqi&�A�n[�����qy�J-#n&܌�@e�v1�&���#�W���1����k�Яj�6��1��KS1��*`�=��gZ�B�H���ؙ@��f�;��2�e�U�y�߀#l��y|g�n//��\'IJ��v�?fu
���+�ҷ�Ƨ�wė8D�"������q��/v� �f@����� on�����A��R
�l�oR�o�0G�-�S���B��!����y�XIm|���<�i��͕4�R����U#m� ۥP��♚6o�R*���è�̆`�M���qބ�/.�����=��Y�x�\K
�>c��������E���p�n]����B�������u�ܗ�������O��Yc/�� H]��}(�F��o%cDW��珿\&-����6R��0�S�2^�鹙�f���&���E�-m t}��N��N�ė5M�؄�Q����_Wl�������N��2��T+}�ڡ.IH~�h�n�/'R�` ����oh�%��Q�L/�Vl�T�h��Q��x�ВG]�.���bLm�^��m�>Y77[�o�V��C¦�3�����'`����m�A B��՚5�(�]��'k'" �p��w��N@MY#�V��%�Ϡ�N��T N�
)�qX_АL��p�>;H�4q�+6���������4V����^3����o�2��4�&���EƸkU���)3$��ӋM�P�~�@���'����\h:lPR����t�]x=qn\!�( �+������@~w�{F��L����t=r��6TH�#D�Fٳjy��͍"L̥�����Ӱ����;n`� ���t�e�+Mޓ� �W3z����\�A~�5�mVW.�l����3w�03��O��������N�DYF��ƕ 5��'�����ڨWx�]�E�Si5��~f0�e�����&fN۸�n'Ћ�9���������z��i������`*�ST��S7厧�Ⱦ�U	t�i||���.*�\~U�65����i��DH�|Y�����׏S���,Ges�ёV΁�?#�H���Mwe]�&�r:�����A��4Q��,kܜF�#�'�y!^a�ѓ.A���l�u �qW1�JS�!��o�'q��ߚԯ�8����:��$���a�����u3c���4x�����M�_�6��Y�?�SY�x�Ϡ�����"��|��-�ʍ1?��k�{�2U�ݛ�ԉNNx����m��\�e��4���T�B��n�:H��W�6�x��W~q�
�Vn�LgF@�:�u)k9�jb�&?�����6N��yip��͙E�Y�J��bʊ¦�~��� ��/��1Z`X�"�F�6�d��,��
�|�fD��Ju��gԂY��UԿ��[4!�J�Y3J�����0⽚r�y��w=��H�quW�[�����~�П||�A�!��LYR�� �0S �D�*�4��+z5}{><kGU8ڗ���H��Qܬ�Ui&� aE[��0TG����J�MB3l�_�2��Z��(5��A� '|�*IP��YnH��h(���F�����,����u�+]3';i���BO��@=xh��>���	6�����1���g�Rt'�}t�S[��i���V0�zEF�ɟ���R,�k�r�%����dY�B��}3���."�;�4h&j./6����R����Ƕd����X���/�>�����$���',�|+�vu�U�gE,u�ƿ��?�����O�p�T�;�)������c�^��v������|68r^i����Gz�tT�l��	�'�7��>ր��D{�.�y��vhy��*����s,/i!��S�Ȓ~/P{ݝ�f��m/�Ww���6�B�z�u���g/ڡO��N�M��θji`�%���j�r� ��sv��k�)MwV��x�,��7�s�;@�5i�^�)�K�|C�# ���{O�r_K��?��0ܿ���^�¥��#��#3r|���EO�c/▹q%���p�1y3�!�_E
���������g�WvB���,�#l>1& �,�de� �Pm�"��h���+i l�3�,��B��3��&�vb��]o�=�'/�o�\4����*TX�y�K��B:ɏ��'ԯ���M&�5��(�U�{�Ŷ��G�rz�|� ���V���4^8:Q{����dչ��b!(�B~�r+������5^*O���~��ɤ�V8g	��n���	R����cy��nM��������^�ϥ/,N��6L/W��U+>�s��Uf�S��\Ƹϯ���ۚ`/?9o�<u�r�.�K��Rf%q�hm�$=��q^�L[=)%K�$���K�|?֟Zu�8�K��kL�C��[T�� H��kS��'Ҋ�K��?�0"�.�w�̾��+S��DN(}~�g���'�H�B����S5
�};�M�������/F$sҎdX�Ed�]F�iQ���sJ����,e��]U��9��;J����]��R�O�D9��{A{EU��y�p)�{��Z	
�(``�� ƽ��O���^�YX0�_N6�QC�LB:%k���\��T� #�%�G��u�4�&���i�VL'q���>2��Ksfkg��>{��[��@��f�������E�JbQ��W�>
��4H��3%���)$D��0�Tt�p�tN�o�%����%MD�a��C���=�A�(7Z�����u��:�"	R<H�Y|Ë�R!����'b4��U��̍ˏN�|�B�˖_��Mp�.C����H8%��&GG��{�3��V��EI��5�q�OV>-[�-)J�d>V��XE�F�V*n��6��+}9��,EL�Tfi�g�3�������y%��y�������0�*�pR�^��<~���ک��9�/B&u�{0mo���K[~�����Z�%�2�C���)��ű�Y��Z�˪�
).���A�F��^��;_ά���:�$L�����E��둯/��{5�E��`X�z�R�@<6��0H��z�k��]q�V�b�J'���n��nU�\��0g,�i�&����Wd�l�V�F-��(�|�뮲���l���	���ݼ;����&1�ġ���n����9�����r�X����#ې%���@�=}���n�:�vD����?H'�/�6G,����p�F�n�F�����N6 �@���_���Z/%\�D��q�y��� �÷���y��5	���F��p�=�Ҷ����U��ϯ8k B�M��G"��H�Ź���3�\;Lw{��6��VW�DR1]u!�*K�;>�[������i���gF�^��LϺ*l�y��B��:����������
J� ��=��H:��'9�Έ���;�u��T��@o�ǂ�A��D-ʝ�B��X��l��X�@��p{��=�̓8$!2D����������3P��<i���Q��8є�4�=�D�A��_|��l:�Vd�� �<v'�z:���x�
,k��6d��fH�:"���	)��z���NtdTc�q�%^��+w4y~�Ԙc$���L��W�����4������b��O��'z�%���8 �x L��]ٴW�]��J�*A��%�����I�U_���fDnŨ��f��.�pˋ�����1V�c	���g��HYY1��io�PT�Q8'
�Bb�Ҳ������M&G���ҧk�"�jmѶ@�����3x�X#��9�b� ��ρXJ��6$�^˟$�N��47uΥ�Ϲ��gP]��ʡ����P�Ŝ�a�߁ ��_���1�Jz;�2���Q�S��ŷ���ߌ�.��r�:����]��d��ż��f�$�sݝ3-]t��ɷ4C:��H�w��1������a�z'�,[�F������_f%%��V���w��!G�^�җ�o{�j��[��_�g��;/n�4���4�j^/+��gN�{FL*��b���W� �_��6�c��1�S���m*^��C�$��6t5�rL��-)��{M��5�{���/`�k�]m=:L�����_��hСlBGLP���w+��C��&w�	@X��$��<r�~E��ޘ��U�����@J�dL@�
� ��VH�q��W�7�nF���5���W~�O�$�#��II������Dˤ��E���AZ8Ǩ�]����V�Sn�&7���X!Bj�VD��f@��+9(i�%f�I�$��M������,��u D"��ñ��ν=PlD�h�u%';H�6�P�wi)�����n�N�~�G��z��wY�d���k��3X�Cw���{��	��@��5�"/w�쯟l{d&�V��
{����~u0'�e�e: SD�QXLۗxkB�X����Q��;��sM���j�G�D��W�'��b��&>��u>��d�bP4���� P&���6���4��IUc��Q�����JV��ý�$)
�n�����n)�sc
NeŦE\fH�g�y�9�G���>e���&�)�],^}E��Y<�V#=�n�_�0�����۫����Ȧ 3��̴���+a�@�#N:�~�%CVIćfBhD�'
�Ô�|�n�΃���.��8����7�ߘ=%�y�qY�ݡ+��C7Y`8��ay$-ר���p\���E�\��ξ�#d��q�������`.(p+�<2��˽�V�!x���k��L��û'�@9^��`����ӽ{;N����:C�y��>,�A*����
�1e��RFPqJ�8O�5��`��$��._����-�S/q����Q<���;B�մk��31��]��� ~uLw;☮����u		U����s�0<��BX�f%�<�G������%&����>W�%T�,B�K�#���3��	�3I3�%�iO�"�`AN�b��1E�(y���=�g��ġ�9���nsTY��H?��Y��ʿpc��YWuDH��]4���i�-A�atQR��#e�-R)ɘ���.V�NՊ�飯�w�x��h����OP��Ec��{���Ԁ���-X����\�,�ݖ�# �ݞ�:�j�a�#!�>J�3�ʃ]�G֒
��a������n�ʾn�E��*���m���\�B����:ݞ7Jr�
�)}�m���<J+�b$��c[�JB����t�^ȌN�.���3���lSZ ���ҵ�~-�C�깯]�ժ��p��������p]����"tJ7N k�,�\,���7�͸����g��C��o[)nѕ�yѰ4/�Y�Io�ai5�dS��6:%i���4ʼc*��m��2;.�4� 㵛�(������k|��{�]/m.Ȁ<��mFB8C����U�	ġ|�:O�]�����̮�����x�����b{�z+���ʲj}#l.�Jl������HM�%�5�0z�ɨ����=Չ��6/���U|X*=&>P��ճ�31?X)����巼.�6pp[*M)�(-z?{&�<_,?� *���q�@?C�#�'C]��T���O1-r�ôD��o'3Z�{h��EIڵjm���%�#�������K�|��GD���!�Z���ZY�%��g\
����&c�{��}/�O�K��}��8�����')mHfns~��&�1Vޟ��:��%�����?�9e5Bz�W6»����k��зd�mk7ca!������D/��^��=,�&�
��t�����̷���y�Y�NrP�b��L��C��(���]��N9��l>��sѕ1�-,�&�Czˏ;�~U���2�?�okۢ�&���Ncܮʛ����x���
mkq���Q)��gp���-s�	����������W��cU*!�h�/�S�;���DsNc ���� �w����̘^[WVtR����w�5�2���jwJ؏+�����C[���ؿ*{�hd��/���+��J�@V����&��Mc�j^�F؂��ß��{�Ȯ(��ͽ�Ц�X{�γ4>�e��on���1^�Z{XPi�/�|�?qϩ��T����+���(�N(����'�
V�{S�d�v�_$ͻ����oq����6��fc�L;��8��T����/,�<[=>4���j�qR�����Y�ƨ�-%����d���m0&�糺]�LE���vv�l�-�ki��*c�4�s�`�1,�ԫ����� �>�ם�"7�D�W�G��]{��*��?#��}с�U�~��2-N7�Q�=/f}�<��$9�p���9//Ĩ�|�PS]X���F�G����k�9��!����@f��ֲ��!i�����������;Cz9�"�񽐲�>�ԥ���v	�,�u��2T�c|�r����U9r1�o��_J;�p���OJ��=�1��q�g�A���R0K[�칎5����1���s�-s�3Q�r�aa���~[U�dg�<|2w>U��m���8��/΋�ñm��.s.S����g��/���sé��SY���TWt�i�3gX�OV��ة����՘�6�h�|�ϭ'6�qR�)�z�#����,���+I�s�z��M�D�;�S�~�^�����|T�f�(쳷��j�x�������i�(r�YIe=���	v^�������#n$�F�sk�ƅ~{׎�7������d��[�ڄ4=��p�`ku�*e��lԋ�jmh��큮��d��:]0��MF�zi��ib�l�5���D)�Hmwm�f�Gn��B�c�{��ws���2�:\,�4����>Bǔ��W�,�B&Lw,E>��>0��9�����z��nHj�g�z?�^�$�¬S�{P�m�ELҬQ�����_������k_�S�W�<����.�3�r�����u�-+O�؞�����L��L������Com���&co���)�`�gq>R:Ye#��o��u��t �VV,� ,�I9���E��$Nn]�Z� �^A��a�l���f���$&\��D�h�"L�\ocTOTr���u���`ɕ2���<����a[QNp����
H����JxZʱ'�|�e�~�m���կ*N�A�6r�p�Z0KW�м�MUg�H1ɥ�n�~�3�c}��!=�rEq�d�d�Kki��3||�IzoPM�}H1c*sVp�i�4i�x�F?����5Ϸ2^��H���"<b��O�MH<���0��Ǽ>�z��Ы��D����3�a�q��B� U��*�iȜ�d�wb���)�Ǝ$��j#�v\_��)�n;Zg���b���}j�'����p?�� �5/ν�T���V4������݈�v_���2�����l�
��E���G��E�|�)�d���
~tr~�<���f8�p���S�j[�Q�����7�
0�B?<�Jxv�;��;��V���u���P��?�tlvƌ�[L蕖&��́�N��63[e1ۛ�� ډUʈZ�qvK�-\q�i8u�v3v+��uՄ��q��~�j��Z�)�����ZM��I���&8N��|�� �v�x=[�){�W]�#N7E�^�^oc�ԏ���w�yv��w����q�D�	D�\�#����?��{�]��k�:�-�}z�P��5�-0��@�eT#�Է��E.�C~kDy{�&�ׇt��K"3�*˨��钦�?�.�x�vD�ˤ&ʅ���f��<���/~�,E�偪k���3A�@z�5�|z�E���:@�i��t[��)1����O#\��~g.K�g0�]\0��)� ��O)��}�����
 (MD���z���7˘4��c�ffC�����#��j���P��Wm�͗�<�-q�iؿ-� Z�xB�еq��L��ڗ�\��N�c�jĩ7�\���y��Kt��E�H��'�}s��'�l��6"_�D���3�?b��i}|#8� �n;�Fr�sR���x#��Ɨ�f�#�I��F-	�e��d������UiUU������+��=YR�}����6�;o����#���e�[(�w���oݶ��
Q�j'�ouK���b�Ә~/幎��_�g�s1��b���J�p)����+*B�ġ͇��'�?�A�@ �N�(�0������a]���R��}�x����1��k���$c��Q?���i�"C�e�ʇ����.����?v�#L<[�P���,b�
 ��P�O%�[]�2N��~>��>��>�ܡv>ힲ �t�
/�H�9+��5%N�^2�3�vu��Ҹd�*�4YH��K����Z���w�ȓm{���{��Y�aa��5ٜ���7�0��R����q�2�i3�h��}�Wi>zB����ӭTV��0�$O;�ܪ�y���*Y����x���>�Tf{�a���D%-*'�[KL��Cs��ܨ~����������v�ND��͚=ɮ�o�𬁢
�*�_c�ׅ_���<PI Ç��;�9Vhjz�76�6'e�p����U�j=U�8�@��X����=>�*Z(�y0x���[�>ܹ�p4�*��`[1Ϻ��oU򄀏�wF��W_L{�"��B(5qUh�&�3�{@��5=ʕt�.��Ӄ.~���~H�
x~a���oy�7-�v�*T�G��T�^�q�-����N�>��ʩ(c����[�E�>��(��"�]�Hwwww�H��H�tw�t.�KJ�s�����?��7��9��3s-�Ar�!�5n#.�d�ɓ�6=�����kJ�2XxNH�{��c�D��dP��*x��@�ڙ���4��8����@m�PCӡ)?sQ�ʐƓgqA������������̴�Y��I	bh��+�2���y��^�9�#ܵI�_�`��@������EI�����w�}�c�'��g.N�7c؄��w���*:H���Wu�<��t�+�߀:��/uB�ٷR�����W'��Ӈ8X�?W���j�^yF�X;�����	ˍ���c�:k���Uo�v��YH/�|X �cC�~���� �74zœ?���ķ�+P��k{��l.+}�}�:3�[����!������L	�����'@Iɭ?�wW��U$}�l�=1}��	j0c��xhp�AM���Iқ�Zzs{���
Du|�="#Y�L� �Z/�����)t����g���{p��e31��D(c[�+\t� T5VLD���5z֥y;�r�k
̃J��
��~��cT�n���s�&Q��F!��"���C�j�@B�L��9_,�h�T|ꌻ���a�N��f�j���W��jiB^�������P4�8�8w>��L�m�W������8�f��Vԁ�t�G~�ກl�����G��7Ѓd�X�G?SK���	��ҶtO28t���Ԋ�Ȏ���½��������FUh�:�=�����ıi���Lh��-lI�+TJ�(���#�C?��bY�z���MnU��)��a�d�}Ldn��z�d�����g�+;�C���9��kJ����\@�y^��c�oX�#��%����Jet��u�M��rk~�d�jXG�*W�Z���Y�����"!s 5�G�!��
`_��"��q����?>�I�H����{�����)(��=�OY�+��Dy�;N�������`�,��2��rS՚U����)6{<�M`��ߩ����v�o���zkG��'u�H�������Vf@�E*�Ǭ�F���B��s�d���ij�[�ּ�Z�c�M���c%�Q�]���ۤ���sܟ�������)Ъ�� t�X	�9�f�i�z��φ�|���{|�w��籱��K_i����zg�֩˃���ƚ�r_c�K�[�f��r6�
�ausm�d�Z�^���=-^��D����V]n�����"Ni����6-��dB�Uf�����O�,C%�Z�a%�� ��� �����*��څ�|�61k����eE�5v�e���q9���Q���/�xG���ݗ����q.�J����UPO���ԯ�?����&d�<�	�Lc~\�3��T����hr{�0^�'��A��~��B�-/��K��2(K
~�ɋ�d� ��Z�CX�wcƖW0�3tT+�!X�L9j�!��>N}5VD�R���Z]	~�?��$�#f��U��n��
�l�j��4T,���F��4� llWs�U���j�O��ID�7Zpfr⻚z��4@eS}({@{%�^�ymt�(`}4���:���H͌������\��n(�8w��@4���	�=W4f���'�TaȦoC{j�<ҧ�W^w/���BB1��аq���Yj���sFB�Ԇ����F+1R�8���������`� r*�ŝS�1R�?a�Cajн*I����4�j+������Cp��D*M�c	�vTl��{v�����񩎟��w�[���Ų�'�pz
����l�!���������m9��Y��q;;\���e^U���E�22�V���~��Û��'r�a#9/�)�;3�Y-$� ��d��Y]74��ΪTTg�-̶�<-/�<0�78@�R*A#_��e�\t�[1tF��}�+�C���&p*���8����JKN���(��plͷ6����}��ڕ9�i���;N�� �5��VS| z+��Va/��+'��[M���[<��I=���ߥx�x=�l}�X�C��;Y��5V@-�JD��<0A���"��Z�=���.��g/|�"��3��r�7�ѷk�� z�H�XUnpU~�'���+��ɔ+k�n��C�I�Ö����.�q'������kw�����U� kk�q}���tҀٜ�/ᡝD�R���d
�
�!�C�%�4��SdF&�o���.C�ߍ���rO�u�0t���3e���JQ�q���f@�*�t���
��������P��}�v����E������R���Z@x��zm���ek:���fʏ.�����d/�f��{�Y�ur�h�7	�!�|�V�&�� �tB���i�rq2͊E�*2��0VEZ,˓��9x���\C�dЏ)���<��w]V�(�yNo�gp�n�s�k��n�n�}��#�e�-����W��8�@\�3R
1��h�oe��g�kA�)�p��H�t��Qs㆑==_p��Q������)ee�p{�^0ۆn��I�a��U��$N��O8��	wa�-È���_��V�[�)����Xܑ|j��N� ��}q��L��t�@�����4Z��8��Bm/�њ�<���,`�V��#��������M��5_hXfO�.���[a���M
��
��W�@6J���Y_� ��n8P&]��y7��"���%�m�������U��]�0Z	BJ[`'��G�:�	9e���I�a��ڌ�8���c�I�3;����״�m��*t��~�>�|E��W����r_��q&q5N{H��ю9~����4�G��?S7��?��BvIQA��σ��ݽ=P>��@n�'֯�����͟
�5����Q�W��ƫsN"s rJ��;dG\�ї�*A<���	ruQ�r�WJ���.E�	�=����4G���)�#ψ�=�t@��Ҝ}�`���r{*�*ù����{�ѵj���h@s�����ٷ��q*�݃�4d�״�����W*��
\q2���ί �����k*Ö0���
���W	Ԭ�h.n��T��Cb��}�(���5'E3��$��?����M�0[������uzAKh�?*�3*��݃t���4���k#��q�qA��vf�;"�o�/�"�Q�	hx���V�$RJ��T	���F�u�ӌ%��| ��J�!�Q
W����t��Jv��ȍt�������2�3g��������G�c�l���ex�����W���p����f,�kݥ#����PO�&�!)7�Q8U�2r��C%�շ����R0�.q���j���G�����Ucr������N�谢66$' �қ]�,O�z�w��u��·y�>����s|u�^�H��a#DQ�sU�e�To]rUO�YТ�����H����tt�����Q'�!{�6A'����A*3ĉƬ�i�C=39��������)4�G��ǻ+[�	�u@ n�2N���8(�p�](���˯yt�e�M3S��Պ�/w6;� ���6%\}�w_�4�mٺ�W�P�fV��'��y ~y0Ewa���=R�q�gW7z������ae��c"ѫw���h�?ƥ�Ϧ��.U� IT#NYh�ɣ--`�������W�:	��(~�E���� �W|"[Z|=X�&]7� �x ue�?��p�H9��e 5p�@ha�)�����\9ΐ��HJ�,힉�B�MsAxyN�϶qw�:��|��p����\pk�
���Fe�ۤo(�	�S �Ɲ�Na1Ki����o�Y�|29�/�kG�W8��|��wq�V���~�����;�K"έ��M[n�:�*�~�aoX��Z����{U$)���1��<E����\�2{qO��Ǚ�&���E�����M����I裯��0 6TH�u�T���00Y>&-���.�P�5��q���R�_�!�i��8��X�$�I�	x:��mDң'0:":��_{�]�`�\�En����Z8j�ۧ&����3���ۀIbc�Վ(O 4$^qi� \B_�E9тk�%�|��S#2����)˳i��d����%<�v�RҖ��it=�NX�D6��<�@t�/NU���at9.$�;�.�pk:�I}c�byV��;K-���k�d:�������~F���cK���@�GȖ�u�����hAJ륿��l���b�}4B�(p2�\��I$O��>�>�b�7
�w7}�o��������1)�D Va4,�@X���Ds��^e(~���l�Z�WMD��� f�]>5��l�hx� 2�`N֩N���?4�خ��I>�Ur�����~�@W�/D�M�t�_���<̶c�ڶ�� i7�U�a�~R�;�u�+O���I���/Z{E��] ��
���1jaL��S�M�&I���g����s�w��C�{����y%x�AΪ<����s��2vp~��4���`��U�;��t���㑷��R	�W��>��g���Q��P��׆t�1���<�ኍ���$#��_�zFx\���T�nZ�3��5̛~d�ʐF�Q!��x�]f���o�����#a!n�2J\G�yy�]�~�&��'�m�%�7��� �P�E�����[𸨈���`xn�����T�_4��q�׍<Mʖ:�7,�ˮ���b���pұ7~�ģ�={��S ����w�l۾��懖���7~��QQ��u�u��@��*e�IK*���Y=�x��꧖��kD[:[�C�K�Z]TX�����@G ��)��X��<Z�&&�x�݀��؏3�3/��r��������E�(7@g|��6�(lrZ�W�@��F W�:R)�!���S�hL^R�/�ѳ2\�=�K1
�Af��dL���DĈL���_�ﮩf�	 �1wS;�N�2��_mQkO;	cwFg:��kܙ�پ��5qZ^o>	�o_��9�K����udT�#	KP���K�ihy	�Zi���Z��������;qF#䨖�~��d��@DA����hd��u��������A�P{�SV"�yl�>��V�1@���k?@���e�q�+C�:Z�Q�S�E ǻ� �vxs� ���x
�	-��l�GʤM}!���F�q��'6���4�����~��)�qql��Vx�OTx\�A��_�J��pS���=3��;N�Z���dZ��Ądh�Z�� ����!��N���J�D�/����<���ܸL�=��#��~i'۰���h)�j�o���p�N<��"���>3�If-���k��g`�O�aq�w�HG�-I�>31KDB��n��@�XE	��o�%�����}-�Wʭ�S�Gvo��`.5�v�o5��|�}jt����N�3�!�ip�nD*� �$n���hn��I���߂��,T��_c����B��Y��� z�b�0>�o䌵v��M�ew8n����Jc+]�����>gG���Qڗ-��p9�Z�&�Ą6�T{�����dC+i���+�]���39ύc�Yy���1�Z�J���^�����ܐ�~|.������wAZ�ҳ�ͫ[��h�/���[4���d�s� �/�/�l~l0���
���T�k+�"�DI�!�����ھ�^�`U��0K]d������e`I�̼�8W�Avi`xOd������^ű�D~c��`��\HV���o�vu8�n���j��X)�y.�JI?x�S� lo��'��,ז&P/��A|m4��u�	�\���T�K��.�:36�B�в��K�v��꺪pW'���Ru��5M�Ζ��c���TtEeVn�O����%�!̛��Ld�	x+9c��R@8D䜨ن�7���/�e�\-8u��<���#ι��q�$x�;|��ydޙ��'�"�2I���6ԫ�Y����EF��5�:X|�ݣd��V%������]�E��a:�R�V�����RUO&Ĥ{�I�Y}�j�K���:��&x��������)ĵ��@ح����ؗ��}Ȅ��U�++����/'���a'�4�d�\��w?ј���~<6Dܱ7�.+��'�]<qAB��3��+5Ԝ�W��< /_�<`���\�Ӈ�!#����򃓍��H�|�}�k�/WeH=�"n�7�6�;W���WL�5	���E�"�N���1�O��h'Q����S� ���AU��BT��+x�ċ�p�o_�3X
O����[
���4�ߐ� �pݸN�N"睎7I�#Fo�y��BA!����O�`�����)������P@�b�s6 f�KqB=ɕ�:D��ē�v��Z��+�ү���F�z�&ݿ�'�y�̃�ٚ���	+´P�D�lv� =ǯ���OR}+3m�V�2V"�_�q�o-f����*���l�dv�X����3��������Y�RWtCP_!��7@���dnٶ��L���5V
r�Z�F}K�7�.*��.���O�Hባ>@I�����	o�E�K#)q�5��ك��n�ůꚨ�$
0�]?���䚖x#�c����6� �<�m�#�/�C�_�Ju�MhE;�;=2{�/�]PR�"< i\�j�wɲ���>�(\�����g	��<��k�p������h*?n0l�\C�6g���w@et��h\^MXD8�م�d�v�k��ۼӹ�֥zgn���+;t��"��q����V�6d\�4�`gtɸs�=����&� ��l��Ҽ��ZpTa�Z��n�A ���ť���W{|�?	�$_W�P�xº�d��p��xo2���cSS_.X��^��g�E�J0\��C�C�_7�osv��s�p�uWrn,O�H	�w�8�T��s����T2�u�*��[z,��v5���}4㞖S�>b;i��^��Z�w_�9��f�����M�{��>9����(8/Ǽ��^G�/I�(�����'єU�7��ʖ4��>��5�?� v-4#���{�Ŭ��]�"�{ :>޸�r��Q4��/�F����̎c�.Zky���XA��[mG�6S�x5�q.C�Kz��W\�t�����[�"�lXף�i��&�_��-'+hM Td~�,e�q�$��{$<��𛺨�>���}`\3x�k���E��}4	��b��叀���^ovd���OL��tӈ��?�$�.B��mP7 �ۭ���ix�VϾ��%�z������^;n�DM�05�}�Hh���	��kG�+O��-���V�!ϖљ��6d��GJi7��u0���"�Ս\)��y���{?Y�e�˷q���4��
NGjv{��t9�p�+�ScFj$Q��Km����{ �I`f��)&F��mӼ��	��|J<���M�mSڕR�@���W�x�n?Զ_�*FJ�xd�~�d1#`�M���+A\�1��Ź�;�5���r�%�S*�'� ��be��%�]��n熆�� ��B"��ᓲ6b���
w<� �i����[$��ߥ���＊KP��I�0Kq��&��?[<�k��}F�}
_�F$�\@Єg廌��vw(T7�	Q�-�ﾭ|�#+w�k	>���e�_�y]jTJ.��[����_�E���CX�?����pC�iJW��.�Pw��i0H���trRT¿;<�-��Ys�vq_կ�K{q@W������L�C�PE����7淋? ���@^�A])A�|ti()(F��9����,[=ܕJ��|���h�r�0���|)
?�v�s���� �@W���}��z�_j�D+�,QĪ����S��%�!��ׄ_ׇ��u��9�m���T\=D��A��P�
tQxG�ԝ����P5�*P�(�1<��o 6)�-$()��j�4�?UVRQ+6�;�#����b��bkdp(��y5#�	�k�u�pn]g
��ŵ��X��U��{{퀿�`J�ʼ���kH� E�߳&���ސ���ȔwXkCCO���bj�x�]H+�~���_v3T����=��95v%��1��U��0 ��O�Ap�t�D~��k����u��=�: ����qf�f�B��:�f�7��F�༏�	$�Щ
Yu�b??a����2�A�f �鋁����J��ͫ"�2��˽�|ߡ��������kÎ ��3�&����ս�����x�u<�v�x�\��[��N�(��]&b��ӵ��m�[�k[�9���2싛���d�թ h�_�BD���G@�)<�>�=�*_��N)%�/�h�4÷f������"�]ģ.��%�?q�p�Eg�%�|�Ħ�8����@�=��6I�;�E?� ���+�����4�T@-�f��2�`���u�o�(���ֲ���<x����{Nֶ�1^�UESj�p���̬�}�� (l��������I:o*F�yj ��NB�A���#�B��Ʉ��%���h�6�G� �$��dq�w S�Ņ<��(h��@�͢}���B=8�����aVv�/�]���E���.^���g�gq�K��ۀ3����=����4%�g���lG{��� h���m�pd׸\FK��9�(C�f�Y.��"�`u��Ʊ Iȴک��ȑ�實�<:ꊅSE���lH.�w@쪍��6�@��T��-M��$���2W�e�G4��SX��<B���6{DWޯ����a^�-]l�Sh�*n��S�
~{�_� �U1�x�������� �(������>�h�qC�����ɺ9���+��U��Bx�~|G�q�p9�O,~>oYe1c��gYcf�x���Prbrr	�ч��Z'�#�@r::�N��%8����	c.q{m�O��VrJ���
�D��$g-�Ӎ����A@���L�������DV�0����?�7�pߗN��p~X���3P
~���M���B[T7������N �F���>g]��u/�& �A�̟`+K^��@�e|�����f�ij�{3���jb42���`CK$�Ü�����M�7wx����Ņ	�ײm��]�x_hIa��c����A�r��X]яߪ� ��+�������L����a�ڇ����B�q_ee��D��/8�����G��%�η��<op2D_�������Vd}��mf�:�X$*Q�������[i\k]E�-��\����Є��_ND�Y�xm ��R���+b��9���\h�U�+��p���}��Ӕ	��6� B>��Jz	��K~�t�'X��L����,��b���_4#�:��&�+n�VyZ���NW���آ�ԋ��=�TV��[$�GO�3��?H��ᮊ�����]�~����|��wuJ�l��ٳ4��� �PD�$Ȁ��]Q�N�:��.�F��mp�6�ƪ��H��*��nq2ј����Â[��bJ��Wn[(�0y��#m��	�_ߨ����C���]M��m2��.�4U� �Jgܟ����k�7Þ���A�m��m�ݑ���g��.(`y���؎6H	�D������b��|xa)Tak$��)���rXއY�������:(�@W�ڸ���h����5���m"C������9�[�_����G=���.͠dZ��Ij%������a����K�A�}�f������@��C���Y-��'z"p�+��T��sՖ��B�w�c�!o����zoE���!?��}�V��v,����&:�dṍT��W�0����}�_�87���#k���s�4�عa�M���]7E]�஍bb�UC8 �3w�� �8&��ą>A��.m&Mz�O��=&��=w�����*T	H�ޭ&F-g�Ç�cT��:y�
�/��J�Ĵ'����j��4�M��݋���hJ�رL�ɠ�Ez�?�mr� �&��RѵY-L����`��r���ʛ��ӻև\�c#�DI��o/�*� Q%<N�(�^c�������D��uY	y�A�S�����u�mȫ��ݹv� ;���8��^�9u�'��?�03�,�����У��8H���3u�kjsڭ�@�Y�vM� �t�vt���9u~�	�
��"��Q����Qj�ɾF��y	�$�_h��6����x���^��'�e�̡k�y���xh_9s�k���޳Oc���W��K҉ ���Q9�� ����	ڝh���Y^�[�s!���+�(��wg�cϿ�T���͆^���h2�v��1
&�mw8��[:�J�O[����"@8��k��>+[��2n�,�/�Ճq��#�&S@�h�<+)+;HA5N�_ru��+�9�&Aü��-Q@���t����H{����� ]T�o�w~�&9�n9���tU����.��m���FQ
�m˼*莯�J;i�Ze(Y @�����+cW]<ksNΌ�g^P���j2UPi�.^�"L���k�*��vps�~CC�[W��_�y�7�2��AJ1fr�/���a�~�3(�Tpm��̬��t����A��S6��|e�=S&Q��XG�.� ��՗+���>���̣�m\�p�ձGҸ`�'���7�9�g����X @ 4jo��_�g33��nD_iWKf �d����ϔՊLxul���ֳ�'�|�G+���̔Έ~\�����N�3�X1�@C��\8�3<\�8�1�/{�I�5tK��{|s�x���ţ�z`I�2O,Ȃ��� W�ɘ�kn�B�U��Դ�����r!�W��>Z��q����G�O�������$*?V���M�ղ2X0]K�s�OL"h"�`"R��g�	>��N14s&{jS)o�dŸ_!b��n%Z���J^u=��msx�}�0��⾒�]�k A2<����k�o�5�CҸ3��%>�ۉ���hP�=L�Q=)\�M`���s> n����5�����"��.�,�����(	� )$	M#��tȆ�e��ӡ�`���<�_�:�N�+*��Y�){@s�`�^>����=�'!
�<��*��Z��竸/��������hў�^_x]�6rJ),jj��y���i�����ک�}��N�N���w@ů�X��A|�-ߥ� >Y;O����e��\{0%٣]�E+3�>���n�xP���Av����Z{Dr��F�Ʌ��)Ǜ,���L��gT���2~_�r��݋��j�<����<5�Snf�Ӥi(�Ŭ�5f]\kp-��͇��'o''�;=�I 9�D4A������e�������A(Ɇ�'.m����_��ݤ��ܩ�5)Ǣ�)i�,�F��Wk��#)A�m����u����XM�K�l�!�[X[[�x��ƕ���q�iÙkYܟ��[U�)�A���H� �N^6);2!@.�:��2W��2����]��=FP���n�pk�W�Bgw�!k�A��I6NO��B��t�%T�������q�ۼ�z9����p:�K2<i���W��}����r9d|3��?P�������}����B�'�!����L���tW2ˉ�YIe�	|�1��{4��ք������`�t�/P�~j'�YCl�6_͙��>�512}z��`2����\�9/��:�����e�p5��n�;���L��ji��-d���!x��o:�OV��̡M
ɴ�����B� U-�?+l����M��L��u��z�g��=�z6p }x��p�)�������R.�𱱶�9�U����A�U���I_I_�AԺ$Z�r�h��|ŦǾ5�\ݒa_nH��n�q���Ж��/�����k�oa.�'��]��,dz�oddyV����/Q"� 3���~��h����� ��p��y�E�b>�L�ӡ6ͻ\��Q10~�S��n4x���"s-� ��-+dgT-��}�|�a�����h ̗�~>��b!�V��eÕ�3��A�/��)O�G7>�y���g�!�g]ܝ��|��P&���;�R�T�v�,��Z���m��C˳ʋQ��	��&\������ֶ�n.��[%B[�&�/dW�?���P �G�/ЎQC	+M�Z�����<�eKkHq+`�;|��U���T�[�|�0�cò?*���lS�}�Y/���l��y���2 o���z3�rk0��-��V;��I���R�L��7y����ב5��/Jx����pV��9��@��Zھ ���۱R����>�ߪ"��sg�P��i��t&R��~�tɧl�R5��w߆.#������	���s�;)F��D
lN�殼5ҕJ ȧ~�P����{�������5m��r��i|#(���:��	� ,I��l�_�H����o��N�U�(� 0���jz�mk1��"wكi�gF����$���&\'��ۦ��()Y�_ںI�_&��YK�=��CJ!n��l��H���K��xG�������t�&D�!�y���w#�HN{!�|�ʊ�8�����Nky��شj��V�*��=p���^���W��V����~��*Ez~y��%Yk"�/�q�:  6�$��(o�����hw��G����xe�)���o�mG�|6q p�	M�w�?�tw�=��W]���c�*�2�F3J�g�D�2�w�Ob���}���G�ܞ��Z}Z� ����~��~��y���-�U֦q4�϶�ش��-L���@G	�xQ�K��%MgC5�Yk�+����� XhFk�^O7Ϳmy���$�F�2�Y��iЋ��zni��lu���@a�iD�W�����ډ �[��	��o���2�H��ѓq��'�Z�$�"�	٪׹s��Ӟ�T�06"��p�.�DA�I�-����挏���Ť���K�BT���K��!��<�O�4W�+����I�6l/�?���qc���C��	2��(b=y f*�q��@���͖iZ��4���q���S�]�cg�H�K)<es����F؁\�^'�Y.`�EG�)��Ĺ	�w��笿At����V2�}�}��li#��kITT���ӥY}*TS␢��*�D2�x��@d��t2K�����z��aQ��s��{r-��_D,�l��	�y�$C/V&K[�}ݡp�����XW�a����g-�җX��L�]�����?	�Z��ҠJB^d؞ˋ��M"�f���EWc��fae��2����S2���Μ���A��_��'곡��z��C@g�#+<�rf����Q �
Ly��1˝�D��P�ڸ��k�6a��e3�S�C)�Y������?E�W���]{�8u%�~a݋7��,:�\����0VQl;�c��ڗ�B)�=�n|@#N�kƢ�=?6�0y�v�c+�]nUfo ��)�z�,��bhl͟%<J�
�\ i��]un�Pb �"p���B���MZI̱w�@���4�u�Vku�.
)��+���s)&fod�r����(�n�z�lvЊ�����zf�0^����ԏ�O�a�}�V�TE��f�t%�ǈ�Ih�%ھîR~�� ,��4���)u����^[��A��ssW�����~ɜ>����!'��ßta*�]G�V�F6��)V?#d⥈ȡF�T���u����������?�3_|�J��S������'u+]�9����y��ɿ|׭�ݖ��:�?��!���X�D�%nߧ�铇·:_��vVP���H 1g]*
�$pV�g=��1ڟ[�Ę�R�sB.B�w]p$}��G��v?�K��NҴ���L��{�	���wi����ۿ��sD�D�7��?z���0���D�pcK�iЩ���ʻ`�؉�~�׎ʁ��م������a+�[?W�V�Iw��Gp���N��0��쪟�Tz�Y�X��������'��8�z
:S��L�	����ьI�S&$]��&�CK�W��$�Yy��������p]r㥴��
�``�Ud��zt�yo����Ɔ���R���vi7�!R�t�Q�	�ҬiQ4;)����-}i�i��e�gc�I����	^��h��8i��U&�jȕ�|}�5ZQ����K(��\C�t�i��پ��}F����F�+�qL��H�F1��_���,�L�]��c�E/�����,��8�(��4d%��C
k�\���`���f��49b�.M&�O�倩d-ا��D�w�yC�&}Z׍u��Y���c��̃�q����6Z%���#l]�u�ꜫ���s���$�9_����k��S帑&ޱ�2�� �N�ҧ�4��G�o~��|�L���["=�j�y�Q݂W..��u�T�P��#�k�B��Gw�Y���'8]y�~����0�W/�h���+P�mN�q��ע{�KW�t`������?���f{��ls�-��
&״�7����f�0��ܢ��IS((Z���s�iQYH1:���Q��1��|�3PG��Q��Z��/�O�)�YF��i�A2p�D�'{����t�����Y��v���*���J�u�zj�&HXb/��!��{��iGd���m�%�'Ō�B�i��h�5��0�0��ҭP�\+^��lVh�\��9�0�d$��ߨ��.�$��w���b�C���/F��t��2|B�%Ĵ�#�/�����mwwd��P�@X�0�S�l�ĝ	�4��%�d��۪:�i��ڔ���k�nSFB���2�sr"#��Ø��H�s���{��F��[���e���~ʿC���[z�˒��Pb�q��c��x�����S�ï�:�^W���'
�q�J��ҩx�g��'��f_�,$*�a�ZQ�����n��L�"N���>�uE䞴?x�Ǣ�&��ڈ8>�2\}�s.{Ü� ߀�`�w���ݰ�����9����T�Q��v[4���*ؤW�2� �`��}'~	����>5�ꭿԅ|���s�E��s׽��d���N�c�#G ������m��q�-ЫX��AG\���/_�!6��2C�?��sS|���ygJA�y�m��+�G\zګ��S�<���\Et�?��ފ'1�M�����XOI�g�d]X����˒��it�Ao�~G�'�·���jg��[����-No.n�<�C�&�]�~$�g��=���$yo�4�L$_p�ϝ׫��^L*�Ol~F���7�����s]�^�,��z�v@�:�>�۲�>��R�f4d�L���An6���w�Bk�K3Vߙ�2����y��G�ĭ� s���Y�Æ�c�Ŧ��0����;6̚����G�|<3J@$r�n�
mT�ދ�}�z	|z�?���(�=��a ����2T��C�l~�Ȉ>2������.S.]�2���\�����>��n���D��a�����L�����%�R��w6t@�����M���G}g��WO�~���P�>�b/@�֬pW�P�%nT��w,��m��ſ-��~���L�q!:�j�u ��tv�����?���߮�I]�q��񦃞.Я㒾���r}㽑��dЮ~�Lx`3m������7Y|,L��6j4��x^'([��F�\�a?(�<�oTwf��*���	��F��o6��ɮ�]�n�e���z�B��/��t��������־���ˀȯe[��l@�v>��,R�������D��bgl]??�Z����tm�Fp�\=?�>?�z��󪞸byEH�&�#�c��0eΝ�8����� #t#á�;W��Ŗۊ�#i ����3//���)ym�7�L1G�f��Fy�o�7�b�sx��	1d�]�3����Z	���c�$ٝ��X�a¿`*�I��q�T5d�:54~r1�p��]ɢWb����V�N��"$�t�p}�=ީZZ�Bh�'t} .��D��ж$b=�)y/0�L�i�[�*�u��ֈ�"Tӽ��b��ZN�1���XNb�aa>)@\XC�3���6�lPY'|[o���B��6��ȁ���wR��}(�/7o�[yDݾ��
�:�/"�'�3�-|^��`�"H�b(0�|��95�
�#�¢�ަ�L�[₧oHO+ޭs=�ENAh����.������j]�"#ꐙ��sv�lG)ԘU��"�鏜��&���A�o��<Z���^���x���+�(�2��O��z��Jȁ"��M�2�gO���
����� �L�tF����h�0�)$������l���0*����.�?�*�ѓޯ�������v��&f����w��f�S�>�0�Z�-�GT�Q#쇟x�{�9%G;p::iV�  Ym�^<�W��jǒ ��o0������.d�h���Q(F����ڐ���a�̵�x�d��R��G� �K�RS2�oj�=()�h߷|�#z~/����T(�NSuW����XFm~a.]a?�w��L�{��˖� ��F���/�9�f4��GoIA�oګ��w���X YtZ���u~B]��:��"J3lp�b�vƯr�G0�Zu�5�����T\n��2x���Ωh/�^��Ic{�'p I@U�F��t����]m���$�iŶ��
0&���k4��P����e��al�$x��w��m��L�4ô�kd�ޣ�����Nf�Zmk̸({.\�YZ�<��p~SN�\^��gc�ɹxF����Ǆq��3X���%zU��j{��g6�/�_�;`O��m���BKj�Wp����빤���A��d{����>�'���VE��9S>{�r������@�� ����5��ӵf#ٻ<�"��cQ��;ceD>#L	���3�L�� ��?�Xp�>��"4�� �%R�5�0(`�ak�G�q���i5�+9[S,U6b{��B�,OC�ǅ%�h�l�^zK�χ��r�Eg���>L}��~Z���(��1��B2�E��V6� �o�@�����.��@�V,ph��3�N�\w	������m�Y���x���vh�놥6�-#��Z�TA���"?��:�h�����>e%V�t���Ȥ ̽�$���ʄ�G؀��������F��������K��EZ@J$��n�.�����A߷�Z��#k�y����o��_'M��r$��!�)�M\缜�Z.v���j?�]��NH	+��Tܬ��T&�gH|�Y�;�(;�n�)Y�ޢ��tU��+��Ҿ�|lUH���H&1Δ���hX&Oo4^�Lq��P>^��<qx'!�NqN�燬����F���.ý� �[\�&d}�����R���B��Qɠ�M0V�}���ؖ{���(5��0�b��|3������ʌ�j�J�\�p�,�wz���H�+g�t���W��e�mY��N<���W���:֥�Y�ur�b��|O��8rR��GM&�4��z��lǃ+�h��ϝ���=b�ֈ�����FETiQ�&����\�Ye�Oߥ��o0�7��^�S)AO2��œT"Wp�G�& eZA�>��Ppmk�pXl���Ge��|�f�$����w�ܺ�����oa5*;�*��ta��� ���a�a��E�u�h�d��4=js�5��0}-_����>޳�J|;�#'i�t�sOa��b@�:���%�d�����W��)A���fy�~�g��|�y���>k���k*>��'�a�e���E)��wҠ�� ���'Hh��Bt �-,�}�2hW�j6W]�p���>@3�����9>���t����j<�^�X�"�+"��� �8d��S̎��ږ�|��\"�Aw�n�mO���z�����6ԍ��ʆUK�X��������Y�<IiJS:��WL����l���-='���b�
Dr�J�u��{�޽����P��\[��������n�����S�Zud���)*}�ŵk̛:�1�^߈��*����o%/�m��p�s]�R�Q�a�o/Ps�_y�Q8��Cv��qm����U���<�ˬ!�dQ�8r"}��^���E`k���9\�����>Q�X��tԌ�|��4u ���[ܶ W�E��QJ�\Ũ��<e�!%0|E��Oq�&�w�DC�ۮz,j��7�D����7�x����~�����x�!ZMHL��|��SA���8:�����8n6���ک��V
����2y��������h�!����&��'m�����;:�-:R�yέ8L \��I�u�e�d���N��.B'�?���,O�?��	1�zc�8��(�?#G@x>���[�5����\du+0�DW�B�l��wL:
;�m˸A������+�h5	p�@��
!^B�15[���[�t�Ł�J����&/B��V����&U _r\���☈���QƀZgg�_
��o@ſ.t��}�#�2�g����H��;� ?1oY/���P��ޓ������`��*�C�)��r�͑w��eFbϑ+�I��p�f���@���S^J�H"��I��or�{\B>+���I��Ms�su<n�]*����
�����F�tɻC�_����?�'�%�G���AK���ʲ\:C�<n݅�v�לɢ�?�Ԙ���s���ۂ��-��r�̞�o��ٻ���q�6��=�O������3z/^���zN^��p��Z�,���Ҍ���Y�RT���<1����Nr��%ҝX�`�"}���M���}-:F�=%Y�[�vʦ�Z�:��V�����?���`ؽ�=	����]u󦮳4��o��Β=F��֞@���K�I����S#������^
(D��������t��%�+	�'���һ�т:���J{��H���̯\WK`��!B����DX9 R��d����������$m���nD����+�m�}�t�y$#���f眽D3��&��ҷ�z����bi1��m��&����.�d��^�����W�1t�Q2)�A����\��"����"i%bx�ۓ�-�,����(p��&�H�ֺn��n)S4#f	�;��U�CJ�F��P�	��B�%,��i��s�����!xԧKǈ}ۃ_�_}���5�^��K (5�!��<��K08�y�iҽ�����Me�h�9�7+�d0j�o	�"t�'����=6!�^�T�o�2���~g�����O����Pb�|�P�8{�C��W�uнk��hz����O�e��Vp% �]��:�=����O�J]���k�H�j�Y��oby�кf�޲��P�n�)��L]˦�Z���CF8m���t�CӢ;w���V@$�~b��I:��w-�B3�����C���i�a7�u�A+��Z4��Q�H�ToE��k�r���vH.J�t��Û��l1��,X6ʢ&
ۆ��ߏ'��R��b>��!�[E��q�d�<lϩ�eܻ�,7[r���dWG�0iI�\�ދ���5�DP ��o`%�vx������x1}Ɵ�%��
�4<�-��C�CAR����`l���ã�{�jyH��+r(v-b@������_��8bY���̻6��-�+ bm���?m.͠�g[��+�1a������<�)�ߎ�.<�%��	����Z�I�������3Ǳ�!�	/�P$/<���:�%&a�_�6U)�!B+g�9^�r5�wZ]��ճ!�l[���ٹ��/�}��3�0.w.+z��'fcuRz�ߣ�5��LUlϚ��U\��*��P8�Z-�]�4���G�o�]����V$J[SO�����zC�U/t�j<~��l�[LkϏ��d���a�,wj��L�Ȍ�%�E�)�W ��M�/R��%Q/
���wG���k�����N�#/G��iN��8(�@fR�"��S�w��/d������V�#�
�)BϨ�r��W]:�+nT�~K"c�Qm��r�E꙾Iw3��\:Ph�¸Kyr>��$"���~���*�FĹL(����~�$����\��ĝ$wPw���FuO������:Mvj�挕0=d�'���e�GhH��ԵDY�_%_����j���/c���%��eo=��L#"E��j��-V�g�b��_K��3��%N�����P��t��Ɖ���Rٖ�j�O*An��0�Wh�f�Fs���ڵ�}�\���r�n`�%�c"��ӰāR�������������?�{/�nxA�L'�&Ô��i-�8�� ǍC[�t;z�9ƍT�(q5��W��޿���<��.ˋ��iA{T�rM `��qnؕ�0嗡���l Y��Jq ���@���+$�ɂ�V����1��s��c|��В(ϰ]'Vp�L������|��ݛ�)o���Ս���Q�n(�y����/��ŏ��L����7�,S.}ޭ�L�z��d�m�/��>'�k��^tپ�N�$�m�ۦ�mc�ӫi�\)T/�<o�\|�FL3�{%>��W`�y�<���T���-�A_�L���z�B�]L�n�?���E�%`��w��\;�a0�l�z���Y������9��ɷ#�v�����P�Iy#R�W~RI��p�^[���9r) Q=�G�><d�=�l���E3���گ2=r~L�fg��V��<BP�B�x�F�匠0��`�*+�/�)g�iC����R�a�[A�fU�j~��E���"�� ]��F󓕫���у��vr�*N���x!�^�0���[:�b��VIvtԐ�S�x�f���3uL�S!�*���ɰ��l����[��~�/�.���2�������<�Q�0=/�\ؗ�|#�M�'�W�S���	P'�m�6���!Q��j��(�	����Kk�N�0C�|�o�
fTtK�ԡ�_���-��ڜ_6�|F��dm^�q��Ujh�,t�h.{4�s�}Կ����9����XE���j�0ckϳ�,�|���3{æ}�P�t˦���R��ZZߠV�5'Gg�T�۞��9O
nS��,�J�s
�>k��}u����9�|���:Cs�|�W���t�n#�^�����M�X&�Y�����Fn��R��A� ��,�1�ާa{���pJ ^���Kk��F��� ���toM	|~�1~�Q��-��Ȱ���x�+Ջ['���\z��sq�����E�\٪������k�sM���h�4K�����S�BIh�+��O�cCv�e2CS���42uĜ?a��$��+�$�m�h�B�z��g6������K�XWQq�^sȅsB��|s��6��fi�^f��52k���'��UT����rsj:w������=btlҐi��Q��=�G�����"*D�q���e�K���KbZY�t�r5���%dRtXԮv�s��Ç:T���CR�Ԯ��������3@�J}���`/ۜ���@^��H'Jq�Hiw���$(��ai:����Y~��v>3����5�⾰�(���������B}��X�tVq��̅*SM��I�]M� f���f���Ք1a�Տ^&欞��Y��1��qz��e�S=���ao`�-⿝�!����T9W���E�܇����/*���Go`/���B��5Db�+ep�J�|�k�]0��{�[CJ�Z�A��T㚭�?�^6e�1:�O��9BH�0^SY��k,����~����V��n�������A���m�����r����`�f�Xߪ�z�o/���6���"D�H�[o�|4��s�V����Z<��ꉳ��z��PV/�9��J�TG��޲�O�X��an��~�l��[� u��W1A>�`W�/����H��|=�t�q��Ԥ��l�"FG����V�"��������q�}�{z�-�t��#챤�W�|_����l�s���T+0
�`].y�����6�NͶ�;+d�<�6�y�)����M�����-o94���r`=潜:�==����\���C#�)C��Ǜ�U�F�-FS����°W3�|b�<�
��fbh�̥�^>�z��v� �Xq����yO*�p�_XKm��߹�(1���Ɗ�ׇ��ґ���)^�A��>�Xx^8I	�@H�>y=/�x>H��z��ޱ�v۪4�(�Wz�ٔ�>��(�Z_؍mL�Ҝ[>} ��=&�ށ|/?}����=�{`/�i5����M���N&���gظ�*�a��j�h�zę4_�vf��d�ƃh`5��KΨ�^��'���dy���rO��P�Ì�❑>�=z���'�za������z��� �4�b5	��ͪ�{QF�{�*��/�D�6��̙�\T���p�g�}8.,����Y�1�/�^�2اX��/9R*Uxʤv]kW%��~$�}���[�/}W7����;��*��>	�+����'T|@��T��������|U���&�M;X�+��6��{� j(�w58��R��(ַ��؇��1����WfL>,ߑU����ﺜhS*����ei�r�9����=|�S`^	�e���,Ӑ@>�+辌����RR���͈"�[b���הH������Z��xfr� ���G�`�y��V��T;��+�i�X�J2����<�����5��k_�?;z��.�u���� �ø1�^��߃�����3��߽�YE�('W�����@����_9k�iqdڈR���$E�ĴAC}�*����ui��j��j��V�L+����~thq����	�|Xo������q�R��"�UlrY�n�M�kF:g�@!��L7�h��_s�����C����S�ʕ�������C��aƚ_M�����1���$n�y�KxR�:�E��SS;��=T79��{}�|Mҁ�,����:��yv�r?|3�������m[qwx+�a��rF��E�g;	L���5�$���v(f7�Ů�s�p�����']��#~r�t�v1���5 D���ާ�f����w��f��mҦ�׭��6�z&9�w��wS*g�q���b�,QQ;��92PGW�0`�8s�;�I1�jgʖ�6��ʂ�ټT�pbs�D�D��@������qf����,�Ʊ���?K��G�)�^Ғ-�\������M�X{%C�r��6'3�ǅ�d�juN������d���n
<^��ȧeǗ�� P�����q�c81�q<s�f���S���1'm�`�1�܊�"�	���TSń� ⾃�`מ����&z�v�����l��$���I�W��k�*����1��@yZΑH���Wia�g?7��{�x����J������[_��6MA"7��M}{�/���A�4�^��=kϰ��bz��z;gO��4��=���#0ëH�����k�]20���_a��D�g��u�
�7���ٙi���Ov�,5��<�@׸���S���U�2���D���ǔ�p��,S��^*f��n�C��Ȃ9w 3�q�M�/��Y�~��Cئ��J�9�4@��
���\���R��$͞��j�Tٯ��6Uv���h�P0�e�K��+��zUV��Kh��ǫ�I1tC�F+x��oҀr�l!�Gv;���2=�"��?GD��	8|���_<��%7x�|�.i��%.�PW���+��_��&�	��tlK�f��P�k���&��%uqɬ��Bwr��ࡕ���X�䅈�W� �N������o'��!W�Q:�=A,L��aG �*~#�,-���#M�Z;�D_��e�s�#
��|��k�Yl�B��|<�͍��?�[��om��JկWz���JT�����1�u��m���8���^+��3�|�^G�g����kM*�~�W�~��y۶Q
"C���[;^��6�3�H"St��E�d���
���ܹ�����8�/�R�n��������O�� r*�\��L��>�z���ZHjf�����ł�d:�/�?~�s���������#�Î޿~��^
���@�g*0��li�"�-�aA�:3�0�Z<v����g�qp�� f(%�#�7]�}��0}���A�k-L_D�Bآ���£Ѭ'�fn����]��:����h�UQ	��F����ż
�����v:xr�,�^_�r%Ī�2��PhÐ�a�QT�C�{ԧ��В�<��B}�r��a����vȌ�%�ͬ�iv�m�hE5#+E�(H{!��/��ص+�pߌ�k��s��d.�ʕ#]��S?"}\�1[�ֶ�=��ʢ/ʜ����&�QD'��&WnX}�x���>��0]�m�< �w��#��	F�;�藘�;�>��mZ�m?q�)������n���L�C�1B	��uN���{�B��� 1:��7���-����{�w`��e��~��X";�$Ə�����7��:�c�M���^dQk�a@V6p��r.�����"�&���_����%d0�:餪w#���\�O�jp��JټBc�y��l/{�(��wӆKpE�3���QbqV��u|)-���ܰ�� �*	n�*ͤ�;��o�� ����e)�JyF/M�U+�>�U�<��D�M[� ��.��4�՚$Ж�FK+@��]�S^�я
��*��ҵ��q���L����7ez�:�!��-(	����/�,���ը�蒍��{��I`7��h:@�r6τ��3P�q�n(t$p��<KL�`/� ��rä�~U/<�DW���Co:8|w���l�b9�D�±�xk�[�)��]�"�	��0�E�?�T����H���?�ڸ��(���Ip������������Fb���$f��B��,+@9�Xڕ���e��Ĵ{(��ϋ�ğ�+�i�s��F�U��g�>���+6l|Xe�TE�׊u&���>�n}H��G�mn����������lY7X�WNEͨ抌3W��^�.Zr�����a��Q��ވ���	�Py�����������"���5]�߉�n2^��hy�F��������i~��!�֦��lS�.}3<��p�;r��Q�-��'��qK�sV��:G-���er5^��s�g�C��j�0�Eg�q���hm���4�]���f���U"[܄w$�c XȄ=쀥Ό��6;b���F��;5nϻZSE/�I(C�쿋�}�Rr�$�~�5�>dv���K2�XN�![=�:кC&�^� ��>f�D�#B_�ǅ)9�&�k5�Y�������Z}W���&��rfW��'�����vP�Cs�󰙄7qL.ю���r���{+^̛9�;N\�1��>����nЋ��� �ے���u��6���#0��{G`����8��]��F��XX/��F�#Y�z���T�"�[�C���T���en祶�!�>�>w!}8�Oͬ�K8��G���5׿PG���0�;ˁ�^��Y��|D��tt� ��I?���7�D���K����_���3 ;#��B� ��ײy���������a�o+��k&e���U�'���Ŕ� � !�6��a��{�V��n�������o�Œ���C;|�$yr��}3��ے��Tp�!Y!�nD�㬼�;u�2��}��6�D�8pz#2`���iXl9?^��Ս�����c�1iGm�MK�Y��+�����P�p��
~r�9��sw�IqQ�`��c8�g��k騏�W��{�/l��w@�x�?� }�B�Qd���dg��w֭:�P�¾M����yX�¹�̗�>�-7��x��G���$�sa*��Dҿ�ߕ�7�ymq��>���O���~���!�Q&� �����׆��,�LoZ�h��}�����m#
N� �)v�����:hn�k��_�z�c��6,��^w~->T���k�3|,��=��k�2�w���u,v��^��a?J�N@���.
|y�H�(��x���1��d�v���	�D]5k�8�r���{-����~ �wJ�/ƍ��P��t>]0^�k�wS�[���4����E��Wj�#��qU���_�3H�)~td����4���<x�_��`ۻ����a���� N�/��a� ��o��>]z(��p3Km���c%�������Wd�ru��3���`��W�J`%�8Z��������d��4u��(�NV �2�q��|Wz�L�TkF ��ğ�.r�����|�y��=�-gǭ+��p�s�'��A#�(����w�y-�2�����̋�u�KGUF�_q�,�]ހ�?|�[��\΍��|����Լ2S���m^9W�0�f7��9+�g�$D��}z�(�E�6�2GB�c����D�KJb��d���{ ��n�}����׿ZL���%��c�3��� �X�*)U���At��u�h6Mh��4��Cs!������I7k��'%��Q��|��Z,�)�}��f+�{������q����nL��~�[���*��P�0ZY�������_����p%�V��x&W�X�P��Fhx�Q�j�6�9�ˀ�R^���>����|>�@�S,����C�'!# ���ފC�Z���y�G��^I��=��j�����#i6�3����g��������&y�����n�t�@e�k����>[6O���c"��Z���tFz�cR�7t��p$�k�	�LK��x�gAO5�����'!����mf��-��bf2�2�w��mȬ��gѻ�i��H�[�
��X��py�ز�rz�v���+5B������P�'q�~-�w���A�s�P*�La�?Ғ-U�-~:L!>���n���	"�D�f$o��2"'V҇@J�� �����)�s�t*��K����l�\GΞ~���˞��D��X��h��G�|�}gw�~��L,��KK��*�Rf��c��;Lbz� 	�"�[���W,����Ȭ��%�_2c���<��!��w}��_!�;s9��![o�4�yXg�O�[ٗ�G�5Χ��OU�zB�������9�+E��>��^e&��f ���+W�ϴ ��ȵ�^��V����J�(�=����'����i��r�q
�i�u���i���ᎊ�ٙQ͜�Ff`O����|s`� ����[����w� �+`کs�}6���!��e���w\�?�C�@j�:���D�ￅ���������ͳl9C�	���/ݐb�{п����w��x��o��:YD�"H&�E�HJ?SMq����D���#�4̿S��H!��
�(C���*H�
W#��?�##�1�TyS�v(�1S��%n�3��y��ߊ�#D0À��I �3��k�k���2�ϵ�����~����󌚨RwP*���}/�U��͈}��DEG�� ��:�*�APejR�?G��O�%ܝ�zU>"Qԅap,�`���s� J�)1i�a!�7��1�%P�=f����^!���x������$�܄״SlX*�qOP'ܛ�7�[A�[5� �Ў-sf�����f"��"hk��=?rb�@9��8���J��=���d��3W�ڙ=�L:{&\�shA��&�#���$���r��G���(���c�V��y�����)Y�P�Q�s�]3�N��'�9�_�6{�>kź�*����gㅗ��J��j���naN� KE�8!��KfkW���*y��:��l�)�����y���y!�'	f��6k�[�c\ys�Y�$��Ap�8|'EH���z� ����#O�&|����q#c̗�� l��<� ^���?���6D��f�$������6yG�Nzگ	�R����@�������i�hE�[*�B����y$Yh���.X�Yp��m{��MV�鷃膱}II�H�-�AH{�V��"S��yw)lo[!o���H��`��� �����u���0K03�
��'�+��%����q����Q��t?�������3�o`?���a��;�`!�>���a��=g=*������ߙ�c�۬��>�Z��}�͵���{�%Oh����lǷU5�����I���g�6��(��Ǐ�L�mjj~��$N����W2���~�#�i�f��+&��ⓐ_�u�Zu��tj�g�R�����]��\Lf���|�\u�;O���2m���/t㩤����-B8���l��r�O��=�� ;Yw��w߉��u|!��nmcZ���E��t�@ő�@cǊfs��?�I_Q&���_���BT�	\+><G8@���9�Q�]���<*w�D�v� ��^�T�#D5-�(�8�\4T�0����k�w
 ���ް��G��Λ��{�=ʬP��z3e�j/�\=���Ĕ��'�q"aҚ��}V@d�c�+��#K�A��\9ۦea] ��I_=4��
�����.$叶�mqN�/8�x&���`x��E6޼�&�ٚ>�0�!�=�/7�P�#P�hD�É��K{���ƅ�d7/�V��5�.ƗS�:�	+���|��Y�c�%Xyɇ��ĳ�d:J�P�0��������ߣ�81����c`Oj�*�W��:�#��>�q=|Jx�Zw^c����N�>
�C}�	�@��[�w�,o\���T�M�IP%zϝqm`��eC��O��MG�WTF�8�'���=m��;ֿ�x�z]����:D�I�/Q@��� �~�@"��TM�DP�4,}�\��zDTw�w�4gC?;�DK�}8P=>H��S7fL�����_L�H�㺗�a�N�q��8ky��s/���(�e/k!v���.��ueЯ��w]Mo5����S����_6<r�eM���~&U�
J@�I@��fw}ĸN���5L-Ť\��c;����5U(p֐4k�	�3�G���:������"PIz�]����\o������N�N�U��yw���q��^M�/�@a��k�e9��@��1Y�zz@�ҁ������	�+�UBj���#ƕ�1y#5"�ѭ$G�mX�Hо*�W)u��(�X�k'�s�2��_��� h�Ј�ʓġs_=���ύ��ЌQ=�|*������[�P���*�+?�q��1g�#������?S�?���7�
�}��^Xx�B����]$IS6�~�~��S�ݪޟ�?��C��N��N_c��f>@
Y���=����s����E9��o/@��wb�A�7��u"��}�j��?�ɹ�+�
HeR�P�~�(5�x��/��<���E����3S��F�&D��0&��G�d��F��S���W��o8�H�ڀ��[�t�;P~9sm�ȫ�F�_�6�jǝ��YW�nB��\F�[�����x�Ᏼ�%�< E�����#y����O�s �v׷��,���ɻRh+Nw��+������Hţc�}�+��i6,�.pE\��]�ݸ6_��q�Z"�W�Bj��W<W����l�����J;R'�,���b�*�����~zQ�Z<�z!��`����L��tI9�@\�h�:�0�4�ѤX����z��A��� �j��Io~#�*�����L�oY�a:��������.�K�� �DO�~����TCƂ����oU��<��-�:B
��v��iZ��Ιd�p����I*~�a0��Z����Փ��`�u6
��m-�������8 ���N@z���l��`��1�	
v�y�8�x����"-y�Tk�,���Bez��Y+%:��v��I�!������Tr���zFl8a5[��t��g{��"�ݹw���_Ú����%s�6C�R�(��lfDc�������>�l>���?�;L[��(x�7xC�w��]↕ܼ?P�E�\����U�02�j����1{��ry���ʝ���M5��涷o�`��A�:�i�l��y���`r�Җz`����62���|?�G���S���r�p����P��l��mb�j��0^�I ^R&���J,'Iy�z:9q�]]?��lph~��Äd��ML����U;�(��E����~���_��%���h:�5P8 �ˤ�@��X���BF�r�Y9}��ghc�o<��f��̠��6
� �}�$���e�Ђ��e�B��K�j��?� x�ƟnğC�>u(�e�b�U�a*����:��l�)Ԛ��Zި]�U�EЬW.��qz�B���!ί�̗:����jo�}��Ca�8���ֽ8u��0%�!�.���hB�n�o����ʱ�>����{�_�Έn7�G��w�r�i��G��$UN������}�#�e:���!�xs����\����e�2���J��"~):�Ď͉Q�����1K_7�lr�odkmy���z+FRa�餵��^?eҭ�!�s��w�֦��\���M��X�Õ�|g\��p���3xSmί]���HFa��l���W?!	ds�D��ꅑd�PeVS�V��3�x���@�Q���џ���[l@�e6%�-�Y�
ж����v�XEn�$S�P�'.�և�iHݦB�ޝw�^�� ���Y��18}�*��W�:2�!�S^m<ش�~SȮJ��5yGm]+�r���Vo�A/ ���"��"徭#��[��I�K���	 ژj��<����kޚ>���E^�?�7$��T��ժL�k�BHʎ�Y���]��-��&�N��E��Hʭ<:�юF.j˫�X���~��g,�*��9]�M��i>��Y#D�޲6�4��n�� �H���� �95��딒��+X"p8/��Ҫ?�QP��e����������ҍ4-����M���)�E�ځ���g���I�PS�L���2I�2�D���'΀�� d���OZˍy)��\���f������ut����TQ�� �-.�ǐ�X_Q�ߴ)��c<���P��jVƸ%?����K3�����B�aqH��'�㔓U ���r�H$�5�^��A[ =3K<�v}:d��_��茙�FlƋ�5;-�>�;�K��J�hIc��Jk��Z��6���*`2��_#��<!/��#�.�����)d[��[�J���pJ�ym�~|�A�tK��);����ýg�qEKG\Jl���p�If��ꤕm\mF�|����Dꢴ����ͼR�{����bb�k��:��_�{���P�̇�� [WZ+'Ơ��?F��h��,�T�˨
������:_�s(��V[F��ȇZ�@��4���!eѪ�,���/�H�X�@}����.��r��V�ہn�GRl� �j�����襦��*���x�ﷃb_:f�'��1�5y����>�6 ?��b8OQr�$��h�ᾪ�ϙ(t�����W+w�,/d�e����%��Z���dZhm8
]��?o�����.0���\9o�c���͔R�����p��7��s�zoq�-�	�Q��.m���̳h����qHsnY�Hv}*�g_��DA����n��C�7_�ZJ�j�7o����X�!�@/\�ry��с��w���<����L�0X��������J\��$:R�и�F�:Qqvb���#�`�l���_�8�X��y�0YD#UiO9w����Z��ݜ�|��Ȁtz��Q�-�x3�n �GwqW(h��]�T�0e��i)r���c����ed��	���gS��l�y���5E�3FV��E�b�[�N]ɇdf���̙š��G��(���`!�GDF��q�z�)B_�)w�̲����;��j4�!ߣ�g`m�G޼�,�n{,d�VjͣM�X�1�44WmP�e�
V�G�xD;Q���ZW˨�۬�w2x{[���ٗ\Ϝ��_�՞ύ0-�5X��Z�ԭh��̘�ןU �'s)�6'�4|�Hw��r�r��t�ǟ~T8��?���w�qX�����&�eR�Ȱ+��I�akZ�
��nэ7�W&�CbG�IƄM���\����+��-%o�k=�΅�|�	����L��mo2�"�(ZM�/�Ӌ!�O�8t���$Y|�/;���:r2����H��1�\C���u�E��L!���/Po�|~���m��B�i_*d�f��-�N�c �J���|u˔��ۦ���V�<�@G��5��&r����<��mq�#��^x_��)I�2����z9	��7�7P,�z�u�yx�t�Q�6�gr�qB=L���% U�,�,���:�:�O���՜_���O$��bK=���M$I�k9i�;0b"���7������?���+�Z��J�6����r�5��w+l<�>_�T��lJn�qn�-}�\��E�G���ƍ��J%�c���H�0RJ��5_�c �WY#<�؀�pg���|Ii���61͸&#��tC����߳�u���g��?�*��mw7���II�/���\���j֯
³����Y�oBP�;��ބ��E2 ,E@�2./��|/t���N��<`�*	b��Ś2z�l��8�$u(�P71u�/Qj�?z�=��Ӭ�����tk �UX�oӁ�����,Ib���P=DF�"Xt��FTuE��`�rt{�K6_�[{��}��iZ	 1�v�|����+=l~�jv����ߔ_	�m��2g���eI����Y
%ӥar�yK��	0���zzh��(2�l��*�	���ĥ���+uأhz���+8���
I�#!�`�$#�_��@�{��y�f�j#P"z�%��OF�SO2M?�y�J������5��N�N�(�ϳ� $�U�X�d�\W��b��P��I}����֔���wl�	�!�f������f:���t����D(Fܰ wW��窬�gs5�,	�^�Z����f���;к�o�[�擇a,��Q=�2�Wc��<��M����;%�	�Y�,���	ލ�O�.���;�΍Kv&J���m<�wN�1E)��̏���J����t)��(e�{tqZ�N*XI�B;�:J��z��± �D����1��K�;p�ƆK��y?���"��'�(�-w�~���lX~�|���Ȓ�e��������(r9 4�d)�Mp���;L���az�&~]�Ҟz�!�������Ggj=���7n�|a&�~بǉ�<38��$�Aǭo\.%��u^iW��JP#?}9`��ԝ�dF�[��6��@�Z3�{\Py9�@�7jX-꫋R��ͅ)��H84�T��������c�-L� ,#?F7��)���T�X�J���"��l�~uj��{�a��D�Ď��fŔ��n@��9Xc��.Ǟ��,��~U>���)�Tр�aSʜkډ���[��=��i� ��.ǧ��A��|W��TI&��-+��+ ��Y�%��U�TT�LЁ�+���x���(������B�2@2��-ǈ��[Bp�N�q͑�������M�Ӂ��/�@��qD�_%�K��T"}
��G���I��ef�j�Xyw}i��nW��A�,mS�o��l��L�o4�qy�Dp	�[��ҭ|���ˁ�'�ߦ�K.�M�?�����WC��!p8�D�9�[�p��!j������]i�7���C�����Y�D<�7���Z� ! �J��ʂ銒��^:��x�&eǚN]��:+/g�{bȶ� �mL#m��}z�o_!����D�/t��*�����s+ˤV���'/&�V�_K�55�ej��H|/[d�Yz{��ǝ�[qv,*#���h6K˗��B3�؆�^���R߿T�[��홳���.���������A>ws$��eW@r������#YPs�u���Un"���y��~��.�>6x�66��4��<�S^��R�!�����f�����F�&��J�k�o�|����9���G�g�c���yΑ	Hf���QH�������K�/���q���M�w��� ����r���Se��@DX�x��aH)�դ��JST+}`ɸ�W�oʪ9�L�:�Mq9a��猴��4@|�Z��[�W���A,��j�.J�����x6��{�X��y�x+�A��-�צ�iVB�ؑ��QC5k[��z��"@�����n׌_P�����stPu�˔�����o(u P%Ĕn�0��nC��D�#����Q>�'�V?�%o���/a�:�JX535��j�ؽ ��y
�=�����j��h�R���t�o���J�P]��}���<)	�[Y@NU�� ߕ5Kz�|�2��O�'O&]};�}�ˏ�����}īE6�,���O�Y *X�o�vx�2��h�O��V|2���%Bշ����``����N9�`#Q ��u�j�Ġ��tDK&M8���T:=)�	J�|X�VcF�^YGʂ_({� d4	�3(e�����$Gʩ��QI��1)yUG�GT�x�� u��9U��e*K���6P�w����C>��Pש��ֹ�4mg�'V��.y�4�L#�� R*<c���g�y��d=G�������m�fږ��Ҭ�B:8E�+�5�ì�G������aQmo���
�������H�P*�%1t(�!C����HÀC��]����0=��3�ts�&�����y�X{��{����؁Q idpw�	z*�O-f�S믷x�N̧��$���G�3��2|6j�z���_	ٛ��O^5�4��R�R��L�s�2�B�������V��d�y/eB���Ǚ��0�j$ ��ar��](�]�}�~]A]6|xz�I��m��?���~گ�ˣ����lbS��i�ʗ0�A�!Rm����<A4��4Pwf�
D�}�_�K^�0h/-�v&���d���[�̉�6�"��B�']��2�����[4U�%�H�u]�GRԵq��A[�H�φ��a�a�^mF��ۏ&����؁iƖ����wo���#7Mҥ�ŕ�;^r�M��0�[�^��ٟf�/�!�(ls�[���o�V�����Y��H�o��.zo}�2	�d��<���ʙrI�^�V��^ۢ�ٌWA�e�i#o�԰Z�ln".�	6Ԓ���hu���˚�$�ԯ������pA�ű�v�t�v~���m`�!,ۊz� N�f������6t~;FK�yH���÷�M�|�Ӌ�b��Y�Ǽ�_�_�)�D�Q`*�^�9�~n��:"ۡ9���z Ù -��I���s�y/n���1�*wt�,��V�q7��(7��S@�GF<~ ���8NV��@Y
�k6�������1�2+��"���MnWj��d�y\��tu}�5�N+�}C4�7.|~�G��i�2��^���)�e��2�%��!�֦�S /B[Hxmw�4z(�K+�!VI��X�;O]�~��4��N����������9Z�ؒ��hni
a����y�r]������B+����49�Ia���`����n&�-��ߞ�ˏQ��H1�tv�A9��/̄*4�ī�R��wT��ր�\ �e1䇾~����͏�5�3&:2�+C��LVYLĞBY�v��=d��Z�_S�z�\��Q^a�� *}��Gy�S5�ꦵ�e��jZ
C]�{��N����M�7jq:,���
v�g[Xn�s��)�h �I��j�.PIb�-G��L����>�Df7�q'�v��.KV������K�#�Z ��,��k7�>�g{K�����$@�P3��e�vuq���<��HF&�^.x��&@K�� �| G�A�-�`��'t�r���)��3�c��9=����:M&<a����ne����'a^KZ�4wFs��p���8���%TA@^�Ҁ&��-8�fG\�I ��
]W�p�V����}<�8a�U�-�w�6Lkƛ�	� ��B���&�]
~�i5'y�!ħ�B�4f� s}�� }�&��ƀ]�|��Z~���7�qZ�o.xF�1woߒ�A��'GH#����
v�r��:��,�A�'�e�?CE֒�����׮���xK�bru�h��T1��a���U����w\�!Y/%lB��\fn�ӂY���N8�QhҲ���9J�n%-��?��k2�W5� ʢ|�#��\Ѽ$�B���̈%��C�xԜV�+]��`x@P��ߊ&���)����C6a��
I^�
����	}�#�B�&��s7�Pn������a�ҩ�O��jn���N���{�B���m`��}�����S{���2��l�!ť�U�U gw��t$���&&A�?"��,���P�2�KAN~d��������֖�T�S�-��)�����#�ՁB<�����ԉ�B��N�a�k�Q�l�2���n��cy����\M�K�(����їB�b����S��Yx���o��IY���y�\��|m�Cl�;�Jæ�&���:��Ws�/�ȝǣ��tBū��1}�o�����@L(0G:Nn���3A�e�)�,1�n�.G2��  ���c.�"��b]��Zo�[��K�¥p���V/��J)e�(�~T���j������rW�,�u.�v���fY�qS��^Ļ�J��V����w�L�w���:g]!�!�d�zcg-�	��ڸRs4!X���ZX�FRy�UT�����s�̭�N ���tY� �:�3�8��F2��������m�x�=�5e�K�gk.�@Bgj=5���c�Ϧ�����d~�Q�\Ϭx��}%1yݔ#��>�e��jp�i�a���^�~�i�{�@��n�]�UPѯ���X���6'�f:\����NL��M�|&�Jt]˾��2</$��s��AH���ڳ������r�O)���@ql���?j �7�i+ii�6b�݈��ޤ���i�f}f���~�UſU>�ŷ�9�yF���] ����h�0�	�NE�s�ګ�L֤��A.M���i�"�x�>u�0����*=�T��N���4������a?(�
� �ycQ���|�^�q#�d�GZ_2#���DA�ƫi,j��	��#��8?l������X��BVY��/�~͉ʿm�������ͺ��m韋���}��<�z���!���Z߹)���^���(���B{����c|��D���_���$�u�`�hG��eD���XwZ�|��4��I�e9����$�M�����F�W���67O ��=�O�=6��Lqu�8��㬈"!�h.��nd��O dO�U-�4�z�}ˑڟX�)�k�D��]��*>Y�َ�J�����G6���aUd#w%����3��+G����e]����u�׳
�{�� 7)j�D.�D+\zטl7ݱ�a#e��=Z(gV��Ί���j!�]	�NG���8)����U9�t/'`O!���D��B�L�J����R�Cf-~�qC��^��5ʌp` ���C�]M�����3�}��5����'C�F+��n�����8���V��p�B�\{�rX[3.�b�$�{L@�!Kyf8C����b#����G��zHW�)��!�m7������Л��-^ޡV^�܁��ߙ��o�s�N��$��ywL�D  ���!HTTs'�����m�f���̂A˫b8�� �g~�\�j��	�Η��̔9t"^�lb�MJ��1��v�P�+���>��bo�:��~&���븍@4R� %�Fe�̌/.agC��^d�g둺*���M.��䣕�4T����6�:e�<O�>r�{�ސh��<���K��ۣ��P���2�-SJ����Z���ʵ��Ri�$��^��^���K��C���"G�,�O`�ˀ��6�g����ܫQ2�c�o�|�s�X�b\<�m���Ya�~]Tg�coo�%z��	��LW"��QP�ȿ=�f��;(ߠ�JF�v�?��
2�/<��_ͬ�F #V�?���s�����C���n8f]��
}����\,R�O���eɯ/e��G�~�2�s����o��'pO��F�����]��"%'�\��P`�K�'����O�����Lhh�� ��R�u�JcB��r��8 ![�g��{�<F+@��r��S�-}ju�~��ZWL���v�fv�Vv��܋�ɻ`C෠�<Ʒ��d7����>��d�;-��NH���ޅ&}�;z ������2�����Q��30K�JEPb��Ml�����~e��٠��/��m�T9��$_��366gJ+��M�7��!��(�꽅&9����O�,�MK��A���_�zˢC�@m��Z�fue�Is��}qң߃Ҭ�H�2�c�5/:{��t��˗38�0V�~|�Y>t/�ƣR��mr�8szm���C�0���w`\]��:t�K���7d� pf�ds��tĝ&������d�7( kݰ��i�J:�}�.�W�+���p B �<�(��}u}j�O���^�U�Y���=�l�����|W,t�K�#�`� C1�E_��B[u�6s.��uN���'/��S�h�0�{#%i��2;
Y%\Ԝ�O��p�x�&���J�ji��	�_��X���X�dU̯{�;Py����	+����,2��VP�Q/@�P4��K�i�C�̡���{���� ���I*�뜆0i��-DQ+��b�4$0���2����t���^��ɔ�Gv(�c��+�3õ �9c��̥1]�+��~f,�4w^�|+%�ꐩV��V"�0��]T�Q�R��o(�<i��6z���� Z�	��B��?������^����1�GOw��϶b���o�ӿ��1�����W��v�o��dO���R��V��]��Lv�$�����˶C�+K/���[W�ZP���c�Ĺr�)�%��\}~�	K�L�޷�/��� Ny֩O��Fٕ3-�T�vSV�i����Y�f��_w�)��*e�����
o�THpg�D?��b
o6dog�\\�e�G��~5�^^�H���P3����,C~��#+��2���������:ɺ���#���"�TF[��)��HP�MP�Q��G�c�P5�]XGe�xFtZ4����R�K�URs�M<���#�_AK�4�Y���Ĭ�,��5���g�}65)�����
�[ϗ���������ul�;
.ɯS m�P��vW��OqL�z��e����!��≯�s~�P���R?<U �/�e��Zݲ+2@�\b��=�����}��xֿ�g�C�/�%Z86?h�9i{2S��BjB��D�=�����J�̱y�J��Nz[p#4��-L�&�����v��sr����6��,�owj�F��c�X��D�?�Y'��.�{�����uc����r���h�΍�U�)D����=�@�.�z���*�#+zMK4�T�b��9����Q�V��By��Mu1��k+dLŴ��X���_E�Od��ǕCy�|�`hbTȧw����N�����@;㻔�3�;�P�e��
��WE� ��w��٦&�V ��鉫9�b�i�h�����--�qG���M�T��r��bZO�Q���fY����n�) ~S����������c��_#�̑��ue@�X1�`8!��mfjЙ����8bAjUW�@L��n����чh�H	��aъ �m��Η��ű[t� ��5]����	�p�oi��0�(>�Y�M>�Ө&�>~�Tǆ���U�~XR��0�A!׏`"�Y����u�Ǧ(��Զ�,���6_�(�ң�>�_ #��L[M�{�U֣�Os��]qͷ�̜�^ϐE9-��.D�+8�b��`[�r�� 5�xB���|�3�|�9��]�}�V��x�-����ŉ�&ɂ��r,��-zѾ�./��di"�L�#�`cg&c�^���w8�=�?�I}6U�&*E��M���C�<Ccm3'��Y����3�a�#��O�󴓀�&�Ԕ@! �dX�|'8mf�[����C�$�Z~��^lu��S�p���O�����n,B�	�)RF l��F��V�4�B�@��wSi�^WL۪��g��&F�_��<>�[i�4Ԙ�R|ͣ��i,��G�]�V�� ��8�#��2���]j(��4장@3Ⱦ��I`w��ˊ�*��z����I�n�^���HF4�W�xU�m���G�N�mH�V��#ˮ�m�7\�N�Z��UZ�堲SQ���o��D6��c%�nS F�!vǹ��W��k��39i	o�O�6����R��H2^�{�1t)$�������{�!^�9��F��~u�*hw���ж7n���"�!��iX���`��f���`���uh��@�����u�j��-՘I��݋�����h��j���puR(�cT���!�|�r�:Q�E����}UX���`�y�{w8�f߈�!���X��2�.K��x×>� �q`ˑ�莱�>��7�N����܈�	���~p������i`�����Z��J��w"I�W�ࡀ�u�EqY��=)����'%%�[��syj���|����X�N���
׫�I����gfN�%Aܐ��� �0Nu�~������U����f[� �}D�eok��2��K�5��g��:lB\?�x�W]f랩{���H]ڪ�k�c^�0~�%Cۥtj�+S� Ͽ# �>0O�%�W�5��6�K<�!p��=�e�M��ʹ6����jn�{���RG%~�ٯv�D��\�x��?܄^��Ǧ���#T@8�!���=�+��VK4��WZ�yRe �R#�����������V�!.�ǽ�	��0D��ec�pC�@K��bƋ|I�	�D�*����[h ��r�z�*!�;Җ:Z#Ӽ�?�F���c��5?�U�{\q����!���;��@~�b9@���*���{qz���$>7�Yxt��'%�9:�&LP�x{�w�Iі�n��ۆ'�VН9%tߤj�=�yϭ�h��������P_=~c8�D>JV|yW�։�����z�`��p�;�k��\�%��>ư����rVݞN�+
�T�ļ�tR�x��և�Ȩ �����%�2��Wc���c�CR 7�hH�|��͢sb���!�>H�s��/Y�'5k�F>��<�{���ދ'���N�^ށ�J�?��9(ޏw¥��0Fڋ� �a-f�?�q�F��t|楓95���{U��>�T/V���c�7��ũݍjY�����3�W�2�� �Ats�&Y�$������ڔ�Iv�NO���L\Sɵ���5⧃O��񉱭�n���]���y�v)T���	�&��y���	8�/u]&>a������3tC�Pc��л��M3v�1��������Q�^���)�K����cܞo���z�f�{�񿮷��N��^�[�~ ��j������ﺇ<ZR��ƨQJ����!��/�W���$�X|uWu܉���h7��+��o# ��6��C�90n��۴>����̲<�צ�����lqf8 
���(3����M�2��w�O:��nf�[�WȢP:9�lT��d~�Z��];�4��H���g .ue|g�r��NC�d�"��r74#7��b��U[�\ݺ�Hw�Q��a�l �@��ۂSȬ='���y�����f~eO�o�x����R����ѧAV���,�ŽuJ��t���e�)��U])f������u�͈W����x�~&��-|�
_�b�L�Ņ�ҡl��Θ��Ǳ���^���6s±����2�����/;�C�2ϛ�w�.tM&�M)UJ��m�ـ�v��F �}n��*(��F��9/��l5&99�3z��gf�nf��
2zkV̜��zIJB�BT�!�N8���*��.�n��'WZ3C ���봛��N(G��m��3K�X�#�P��_�<v&~S��G�hD��|�i�F[X]	-yqz�\jȣ7�p�b�zg��(�gA�K�u%�F�:g�QjϞ�<�����{�kh�VZ:���{\~��e�27݋�;�|�#;��Y!YA?�M��=Ų��I��!���������f_��!0�7�Wk��|z��lPh�_����+T�i��
�����ƢZ̩5.ɿ���z�r��G㖠�Q��W`�`��9O��w�_���]�R�UwKF��ɢ��	C��b�����ː�X%�W�bʉ,
_����o͈�
rg6�}8��������}͊��e�fH�H3
:7|3>V�4>���YW��i�5?;2��J*�&~BC�5�н����%�k1J~�9:Y$�8��Rʾ�j�B�'7�f�?F�狚w��)�|1�x[����^�y�hN����}h��U�D��1�,�j�T����{�v@�0y���R�7��P�w7~���o����f��  Qu�ˋ�����2��G���I�	A�wt�#�U�B�6��\��w	�^d>�M����n�����я[?�3�˖�Q��ne�Ǜծ��P�R��K��F��[�M!�{�sY�B/K�G\s�եj�LʄYѳcY$����yC�G�������(�>q���(�ݩ�6��� d�~˞'��T3g�m�N�dP�����z[�G�Yxk*�x�̚�ɡ����S���G��V�l)�o����aދ�	Ix̀�=g\
@$Nh���t:�� ��q���l�����I'��.>�3RIc�t�c_���5�u�����Sf�ben��Bǔ?�"����ٖ�[�mv�x]}�T���P�~�i� �G�u���]</�υӦ�����
���^q>��ƪ�}���Q�)е���L��-�����)��%�M�͈��Y@(���B��3��d����)F�H� �g${���'s���`"z�����v���߾��M�{VKud�>͈ ���y�.Kq�COE1t�'.���Y�:���ʪ��2u��ZJ�랛 l��HhU�_yZ}{aV)�QS��%L:l��}� <G�*�P�Ua���S�'��(o�uu��f�i�V�� �mo5�b��f/��Z�ރ�p��Vwk�1�?����az��08�E����g
v�*�ܤt�L�V2�¨�pǴ�d?-����-�F<� o�j ���V�6g��mP�x7�J����V�Ek��d��hN��*�8��
��^8~���@H�s��ש�b��9>z@�CL5�^����W�~!���^��7`Πl)s�#�Dl�7��P�&TC�5������Ik���\�4��|Z��{%�zϹI�4U�/W������}(��p�__����rfW^}��k����m��*M�ӻ�����ף���a��E豞��D����q#8�h��Z�ء�Be"h���N4|H2���<��n�Ѣ�uW���0���GS�
��yA�`Cs3�!��X�h@Y����ў84�=����P
9���ʃ!�%�ҺF1��$z<����LT���b1�Ai�ww��)L^;���-�}RQ��6��gU�c�i�;����'A��v|�����a���^=Cg��i_C(�@�%xp�7�S�D����З�W<�N�R+)֬J�q2t�S|-9 �m�r54��RS���a�m�	�*�/ � ��:9s���&?m`��W��5z)�{�`���۾�U��;*�L�~��u�?�U�D�{���F�;���
��@�b���Ǒ�)�)�.��?�ԓc����U�c Y�@Y�!~�4Im� ĵJRD�u�;g� Z����e�~W�1�b��e4�y��P��F!_�g��]y��B��	�}�A��:��UV={s:�&�i5;����Ƿ�՚��3��KGpl�kT.fD�^I��s�4O�~�TMjݲ�T֩�fU{{�Cy��s���#��H��m���e�#a���Y�B�)gK,�
}�3�-i:s��?�Z�)���$]���T����0�It-�`gKY�G�y�'���o�8�WU����u��	���,{����}�R�
��+8����祖`��fbD�&Qj^'�0��O�$��V�wr�t�γ�>��<|���ҵ����&S� ��bBcT������P��c��Ϩƛ����yف쁰��g��S�����~�N3+�"c�U`e��X�T��ZP����!i+���F��3�����i<~�ú�f���
��f�������w�=�g̇/����9�����.�)��
F/j&CS	 ̀���*3e�����әF	F����'�4C}��e�-+q[�%ko���~T Q�d#����|�@g*� -m0����&�&L���'\hGƍ+>�6D�_��Rי���W��rnm�O�i��v�q`��}�.�f���#��/m�x��p$ɫOǛn6�ě��o��sRvk+�=���gUQA4�^����9��ʶ�^i�^�ɗ-�\�h$(������-�`��"����~���L�.�!f~�Z�"v}}X?(�<�Q_O��)�\���ݲy&,�Cb��gߵ���vwݗ��S�����wl�;q?P�;+��((ʘW�B��x8�Qg��*���y�s�� ��3#���#���g��T+��9��Ļ� a+�w�!_�B�đ������]2�W�[�)ٱ��3~�w�V���s.np[dX��9���s��k�ЛdT�/�i�t�垱�2�����b[�)�I���y�aO�]��'o�w���ν�3�U�P'
k���1>�T��I��$�kt7�5qD�9T_��"{���S��)�OΝ�;�(����Q�$����zr�i?sG�!����k�1&�#Bb��t2���n�NF�笖qs]~3d0���Ob�XFB��s)�?��0]�V�w���2��b�Xv\�z��fl_�vyxB�����uF�d-���e�߃��~F�R>ۑ8��-}>^��x�� a�3�K!>�n���l��>�?�������uwy-䑢�T7���5�-�����x㧲�Ũ�a>���l��QC��R]Ԏks��bSS|�%�;� ~�`5Q��ڀ8MF���+ȟ(���k�J�q�_���P7�ӫ8�@�*R}���Q��aɝ��!��]�,i6O>�*Vp�V��3�x�i����^Μ围�.�P��	Q^�o!V�=����yJ[�pL��_�<���\�:�Uq��0��t[7@6�!��ӧ^a���8���\��d�i���J��E3��x3��R@��fwѴ%x���e�MĢ�ZDD��IxaB�G_Yڤ� :}�e�:����k{�x��g%x����>
Y�����+Q�;��|�����';���)��=r�'����`����y
��E�/�Ҹ˩J�2%�vIUe�l��ݙ�ՙu�7,F��p���,z.�	@&�
]>�C���Y�>_��_�����j�9�TDB2�7X��܊�[<�Ә~�����6~�A�bﺇ�jW>�B��wY��f��ήoU�E>��~$O�.����������Vm� �ꥼT�Y������`�O�3=��?u�9Ҍ�q��3�#�W����B�q,'x��#�Z�	��r+0���ɣY��nzR&X�"/޻�J�?s���%'To��yI��GOG�4�e��5�>U�I�8-/��L�d[4G���|��S�8A�Cl4��2��?8[��z�.�dk<��\q�{+D|�Q��F3�v��ؾy|9�z�\"d�n=穦��}y���/=�w�VM~�bQ`=^ �g� x�[!&9���]d����x�1�k;���Ǚ�fԥ�h{o|�����Y�Jc�/�9[Ѳn��O�k?��x��������V�&ݖp���-�+��3���8q�{*�3;�$�M�,��-��BH�P	/�Ԩ�����+�@����Z���H�s�y�b���t����kް��#��=�.�)�.��s���Jq"�o���z}*J�����ɴ�r�����g��DL�կ���<
v1��G���(4�J�7~�6�Uᱫm�DV�=�AoN���Y�	��ҳ��s��ci��+g�6�����Ta�t�xU��e���T��S@�֓�a��8AhN{����d|�sᆎ�.C{U5����E�
�w��,	���wl(ޭ�N�۾#����	NhҡT�c�����S���/īd���'K�<ݕbA#0̶�Iȁ�<w��A���6����. �'x����}*��?ӕ8�����b.���
�Vwv�2sH|vɼد�y{�pp��c_�_�L��i���qY������-������lޤ�L���7�0鉳	� ~�дl�f�y���v��A���-k�B3h�7T'�}�+���9�^���gH,7n0+��O.�����u��(5/�� ~�g�#���3onz�p�}����;U�^/��:mHO9��� c߰J�A�"1:p�Mɷ��c����7�����k�������q-
_!��L�&&�,e,����� <8��KjCݕ���t����h\���4/��k�R۪��v��(�����ȗ�ڴ;0��V��b��!�\b�^�}y�m�W�oQ�B~����C����r����st��*7����6, \R���)��c6#�ރhʢCC�����GǴ�csE�=f�g�k��x���z��+ռٝ\:�������3$���a���P�k�)txZw�g]?2	��3m���>(�=�K��VtZ?Na��Ȳ�(�\�,��{V��) ��?g�9˦L�b��w[T~���*KI��;����/&�� ��5���=֯0yI�G�rENG@e0���Z,�`������	�ힵ�*��Z� ���8{���I���ٸ�myNm�HCo�^&��ħ�S>|��V�X�]�WQ��*��Sz�/je���U3XG]���6��3ξ�zh����X�):���egN�݂�`�*P6K'뼼]�ojj�G���5�*ϰ�G����i-��ʧ�w��ۂP�}���K�To�0Y�*���<��1s����(�'�Ε���j�r����x�y{��|�P�{�)���W��?��U���c������ک��'s��O�_�p���-挙Q�����8�Ib��J��)�e�߭���!�WS��$����*����0m2�N��o�`7l�`����⸘�������Ni�������+1J��vk*��̼�͏V�K��m�������b����L��u�Y�* ���h�X;_9�l&,��U���%��Ηm`,����ո�y�!�9�p�O�̬��J.`����sX	f��7P�F%e���՞��?n�*���ˍH��/e��a{�W70�4���y"j��c�j�*�������&S��*��l�NOg���~�����@L�Z���>cMU~�{�~a�2d~8�
Ux�n>O>I�<����<�:V=;�s��N� �M��6��ױ.�uF<H��n��ǯ�;?|���T�P!�[��g�nh������n�����[�sc"������;*W���w��/њ�ꦒ$XSb0��7W�,A�Rh�jr�>�f(PssH�#<�n�s�M�ۆ%F���P�p�^[*p.��Y�f�|�Yǲ7���w#�H�e�CaŪg(�A��X޼���r���n,�n����7փ?3 �R{�t]�.*�kY�Q^��o~+�5���O=��2o����x+;���}�j����bb�s��\�lw"g��{�y�h�=o`��I˫ę+��N�rܽ�$qp�D���+`o�Ϥ,T��_K,�Q[��&�Zhk��L����,$YC����q�}>�j
i4���ܝ����duT�he�T��rM_5���XG��U�k�-2��W� ���)�fę�j������� ��
Y��<�������@��4����9�֗��W�_��K�>u8�'�3������K ���ف����9�r@��9X&ӴT�Z¹F1-�r��*#{�t���~��>�7�^�]X��}�^�ft��v�
�� Qܹ)��5���p&T���uY�9oE��a�Z@VB��"U.�)Ǒv���ږ2��!+-�^DS"dvIӌ�O�� �ӛ��xš\�z���Tl+[���\)��S�|<X��&M���1P��C�W�oH|�Kq�?�˨S�T�gWL�Iv���K��~���!��#`�#9��ڣ��U���W�ߞ@}�
 �'�95�/RT1-�T?ɠ�PLo��r�$�ݮ����x��K��o��A�
r���/v�&[�]{��ej��"3��8����x�Zo�ᔹ�ݝ����wǷ*u�7�I��F%��@�2z��dؑ4c��͊C\ ���E��6FG�M�y��R/u�o6��pה	�w�,�����<�@R91\5����ũa�җ�T�}pwTrBP��1�0	K�N���=y�!>����X_�a���������_���D�7�ݮp�P[�*C�@I�?/�Hx̲\[�E�$N���#O��_|���}���=�R��y�xU�Pj��Kl��ȷ�nc|�]kpl�:u�y$xu�X�mw!�S@�qj�n�,�ې бa�z��׮�%��3�����a�/׍>D�������+�o�<;z��ߜ���Q�L�/Qj�8'���D�K�kpT�� .�Q;���䘦��ò������)��C	_�(��ٸT��:��`���D҂E��_���гT�2�MI���B�m{T
M_|׺�������\|X�K�J�����Kfu�ҍ�3X��]�ft�@�����w�ߟ2��u~��*�
,.p�qM��愾&!`�F�� ܢ���t@>�s��/D�{�Fv�E�v��n�8!�tͪX�!!��&M^����L�8W<�pI�#��bi6��
Qh�B-�X�k2T��3�'�Q����$8F]y(�ۀ�1H1ͭ3���o�!�:�%X���Μ�+F�O.��*g����Oe����0�T��0�xM- A�5hk$��� ~�Q/>��e�2*�k ��[��(�����03TW��m��4�C���Q
]PNN}gO�$��q%�(�!B�X�$\n�y^���`�m!��	�Cy��?5N@Xn��$�� p�
�k��7O�I7�*fz|f`�?!h�}�p��N���J�(e�qTڳ�J���Y��DH��@�(K�����^1>20d����R��*�̱j' �rJw�c�X���!��\�<���Y��h^΄tm�0�[5�
�楗��ۃ�EoD�����֮�hcL\bv��殤���2�Ju���Y=��y ;�p��Nr�jMu��>u�g�Ie~��4�T��#�S�L�3G��os��)���:�}ew``f�u3@���kbU���-�(�m����v:�s�;'�
�K�p��v-��.^�G�݊����Fc��S��������(���yL'��oGX[Z�W�|t�B���ռ$2��5<�GW�S';����϶ū���'f�Z���J�ιI9_�,���fP��GH�s��9U��t����e� Zd�$VT,]����j�t��*�J�5�w�QE rԑ�k]��BX�K�vf����[%�W�9[?%|�>�B��!��q"���.g0B�qJ&98�s2]L=�O��(�i���=q�~W0��������6�����'vǻ����cz% �RZ�k�;��M�FU�P:�8V_�nj,o��w!&(����6�l�����IFˍ�8g�&S�u����ƴ$au]�E`���%��o�p�GU���H�m5�lz<�B���@�uJW5�i�┎_�Tbl�����]@r���Ϭ�����F?���׆Yo����N59Y��\��w�[��(�2O�Tx�_ơ̈̄��$&�ь&���ONZ�O�/mpC�:)�Y�Y�=&�ה�OҌ��:��ڍ]|h�1��)=E��ӳ�俇uf@��*�H�
0���(���D�A���I��cɬ�P�䊮W �	q�,OxVH����;��o�o�7it�y;ߙ1���mZܷ�D;�0��"%ǫ�U�&,�W� Bм��6*�3k�6������2�	�ɒ����٪�C��+���$�(�<:�oAm��I��8~#vG?=Fu<tzK�yP؟����Z�&҆F�RsX�ICf:��MOj�����Go�.�y�Mq�4D�x ���d�$<�vrGT6��X�:01UbY�=L��Dx�tCf�1��xĲ.ˌ�Vl=�`Um����?rw��(��vE��d�Lk�J1�A��pcbi�;�lّ����W�؁7��7��e�������7�~�k�_�t�����Oy��%��"���}Ph�k��T������F>;��M����נ^0"ȟ2�`ŗN�syW�&ho%hL�L�-�U��HUa>>n�D�LT6x�E�k�ߔ��3~�U~1C�`�� `�����;��j~yHl;L)�5R��o��"���˵��!!-G��{,,��y��颫�0N�j��sܾ�s���5�V������"�~����ԙ�,�Q(��J�$��G�ޕ5�h�驜�)r�1r�ؔ�pu�-���l�)G���䭺[Mv�1J[j�`t~r��#3�C:��w�g�>�۟��Lb�O�=��R#���`.��Ӯ�tN�EB�
'KV1F��5~��I$��z'�^��Y��	�x�"��y��"o%��Nn���#"����A�?fQ��c��eg�>���iV���?����.?�2�����TFV�-�T4�J-��	<���^i#	}�Q���_ڑCN������Xtj&�l\ƫsR�8Hn���_�l�罐�O�ήdψ�_��S5_���[�h��Z�ƹ��D�ц���zi����$��0q��'�W���P\�(�JE��N�������>���D��Bi!F^�>�h�/F�V&e�63C{f���ҁc��C�Y����?z���<LE�V}�����ap`���VŋtT����"]�#�U,��SGM�$r#J��KwM���4Ę���%Z�a^V1,���������K���bM�lq�OX�v�����_�↷�2��	����ρ1aؘ������'��9j�o_q�o�h�>ۑ��_�G�t����w$��ͧj��9����yf���6k-�h2��L�`��E�·nppK�kze�VyN�0�����	DrּE'�,Y��s����=V�n#wd�tH��ו��(���Ω}��S~����_���̴�@�"�[��+�}�R�D )��y@�u��؅\�*�WP��Z����߯l���wJ�lG��&4$[�!X��XR�"E�������L��H-��u����,��-���߃@�0&�9T؎8��������A���!Ln�Bd�0}�S/�4�8�N�&�AaX�P7Ű��U=�"�o���5��Y?��7�!;�Hi9�g��i�t�9/���:�0�Y�N�%��dy��rnlu�Bs��o����~�CXq��(�"��@�q��#j4t4��'��چ7�&$��ՈU:"�\&w���}���С܆�=N$l䜣�px�d�)�L]����W���F����ފ��P�D��������O�	���U��@"�>O�J�zL���v�KP�へ�� "�����}Y~f����g��U���G')���g�N]���E�M�\�"͵��c�G�CZk�"�_�B-��IJ�Z�0���G�<�"P���?��8Fi>z�K^�b�ˎ�����$(�2#��v�qlkt��_sy;V�-��Ɯ, �Ǌ�,���?�Uَ֋��w��;�,�Q����7�uQ�	�������iM���˓m;Q]؉S��*�ˣ��~������h%���"ʳ��5�C�V�Lv>�{.�P�#����I�0�[;:��Y�w�H�b�ch�ZeN�\�D&��Ip�ì ��4qh��I�G40�_�D�'*G�d��r��K ��S�]�T����d�� ������Y"���5�.>Vr�م��u���pN��j>2�"��ʷ8����-ذ�V�1���Bw��(�rN��Ok����d�[��� ��f�gSr۰Bw�Wo=Lg�
1���X�eP� a�=���a����!{����K��Hq��@P�-�c�YI�0�R���/�N��dG��HՊ�kcs�C���j!�V��H�-�v�?�?�5���e��8��e9���k�������AE&���1���74 6>�q4��8P�5��Ϡ#\�b��Zz-~v�#��� ��Ԫ�x�w0+V�O��u��@b����:��^���f���H�AUԈ�n�����R�[���v�]m!	<|?i�ew���$���SG�i��n���:�s6-%F�Y����.���
��/�`�	�8l����*����>�g��l2IasB�p����9iƿ=���������)K�E�-��f����.��_�XgB�LeZ00�^�����n�cf�48Xr)���E���}ݚ�\��?L}u\T��5��� � �%RCIKw7J7�RR��#0 C7����tI�t�Π������9�9;�^k�=�L�Y�¿����V^V�����T�&�'�*�-��g�j�}G��0tr�_4�����?�gM� ��7�9�ρt�صڮ��w�>*;��I�p��Ac0�E�p��7��ɐ��i����o`��E #�ƥ+삾�u b+o�2�v�����i�(}��z!�`���n�V�))����A�cl��1b�!���;��[kVЁ@��
\_�t�s*��,� Xo�T�6�X���9o�U]�gt����[j�����l۩��F���h��^�b��x�����HӴ8���H�(,�f���(� 8�1q�UBO-�S�O9�g;��F�a+��-�4�VTy��b.A���{��j����Y �b����������U�	�0Ɓ�n�e��s�8��)��C�U�l~�SQf�XuWU���r]�����F�TO#aU����Uۿ%NӞ�5&b@e�����y�۲M�L5����yY��7�������6�z�7l��	�n��ۮ���q	�)�I="S�7�C�Z����˸C���K��bi���۱ܥp ٺ��Q�Ք�~�ϽA�����2���L�B��]WǛ�ؾ�955����|�_�HO��8���/ɱA2B�z�ed�c���m�[j9Q�X�ۀ(A��w� "�S�ۜ�5m��A�y�T�G;�L�M��8~Y|Xn2h5՟���߫�8�nr�2�V~F�� tt7yt��讎�y�sc�>0!sa��f8�G���[͂A{�!�N��v͢��Ϣ_͈3��'@��a�`м�SR��/�[���=� #x�h��}�``��Q����<^��H��C��
C�*ejDE�Js����0�-��Kv�����^̃T���K��Ş�Aw�]�]�hR��]�R;C�v��c�赳�����V)�)-5��:v����e�r ���-@U���@z,�ic<��p|�ʿx7��utX���(�S���Ӥ��L�������&̍�(u��"�c�&13������J��˫E�˫��ur �O��������L��PR-��Qx>�N�����ڃǙ��;�ʙ�p�ʕ��l�Sy4Tqq���UV	(6U��+G�j����%L�+��K����m�x�,���)p�*�qw�;	��v+D(�i�/�H$o���a�£����[�����!ȭO#J�gNG;R�:�G���Mu70��}�0��� A����y��=��6n�|�0/fTIv�qtt]H��<?{����;J��k��qh�ڣp<��k�s;���j��i8�R�Vc�TۥD�l2�9�R�yؚ����B�:~d&}�K@���$P����d��?�D�m`��)�SRkJ��(��K�G.r+B&��U��vKkkϬ1�}2�S�l���؄qr�A8]�U�MX��6�3r��^TC#�K�@�;�!w��JF�զR�N�7�_��摜h�e��2���b�
!yw~|��!;��s��F��N9�O����!j
,)A�3�L  �DDŖ)7�M���#"�ꛍ]}$��6ͳ����3$��zSTa>���1e]� ��ɳ�����E�"��9�� \%ȱ#���|���.O�k~ވ͗��3O�H޾�2���р���d� dn;��q ���R!�;�sjW�`�X!��cm�"eo$9�O��Q�{�[4����ԣk����� o������#���G�d�~���~;
&C��Y<�!�����&�m"���&�@b�k��X�����	��A��^0����g+���]�7^̙C�o���P���)�n����[
���V�s����f��:��{1�����~�l��:%N����f�F���FڣYM�!�{g(����hg1DT�'1]��'�c0	ᦖ5a崻��gD����i����d'niU�5��Z�(�o�!�X�|ac�7rJq�������w>E"��g�,��Z\/tb6i��� r�k�H�Nn���B�{��X�&)1Ͽ�0 ןN콩�oT�����>����q�0�d����hO��fxM"
Gb��$�����ʲ�>ql��_�8����%���sF^�d�߂ET�?:~]1��:�k��.������z�٨��c�Sr*4����L�-ݨ0Hw5P|��VY�
&B�bv!$���6�(���٦��?�J���XU۽ڞ�/�Vh�E����ǪGA^�2&�$3������R�""5���p�ւ[�M�����3�X�i���s�" �a'�G���a,.�!g��u�<�b�9�^�U5�kLa�<@�`+�n(�)�*�!���?�;9������p����p��	m2�1D1@j��`���F�	I�n���<��/�y�H{�U�6:���FD�x��6Kl�n�?��Zi�z=��t_�\��!x���~1"��>�,|*�x4�68	��� ��� �3�J� x��^|���g=շ�d������g�͂�@�f��N�� ��X|��\���" ����;�Ly��}����-zl<5,�pH���f=v��Pm�_�wuf���$��S�7pD4��"{K���I��.YV-�s|��߱#�iW�#��Y$��~��>�{��I*b+��AѲZ6���2�]�f�[��X�;�y7l��x1ŧ�\�������	ȕ[��O'f��y28SE_�ˌ?xBDr�y�m'�K�=��oe�i�|eJPZ��9>��B���T���O}�����X�&E��(�M����J#�wG�AL����]��!�g �y~_��[}�oa���x�6so2@<2_@�� 	r�=��~|"b~�����ҩ̌N��k:@�!��kf��f�i���t}�Q�A�(���h����u�b!�o_.�5Tm�X��\�Q!~Ws=�g�v�fGզ���̢�6���Nfs�� �I0���̻�4��?O��XRG��2O��gU�u�QRYћ�-�ן5*����efv��c���:x��p�i�1#�i]���g���N�����jJ|��:W��e�M��9~U�ED���dHvm�I��+�X�E�J 
5��3
f��J4�����^	�J�-��%��� z���k�~��:�eo�9z@)`����������U�������b��%�*ULgV�F���B�g�@m��(f��@����~���a �i+���~�{%��c�O�`��){�����A�L��G�خ6aΊ�������z�Ӗ*��G�H�� �8���7���4�8ſ3�>�0�%��j�]�8�N�[rȮD�G�1����\��S�{�V�+s�L��TwŨ0 �3*;/,~q� �d�p�3�s�������:~�b�mAf������[	�Z!"�J^�(�Z�4���C��abz��?��*Z+*��C���LV��X<*�AL] �H������H��Ub�.�wBhj0k�̏���N�heC_�q��n-��F�;�N��e���c��ƗKz��Kq�`����o�eQh�ӡ!�[������l�l��
�c�����<���6�^��I��l�1��u>Cm\ֈ����~�(%$��5q)� �+[#f{J65�h���Ds�|�וV���B�b��@�P?�Z�_~�_ ݗH��l\��!�/#O��˝�5���s�ۍ�Z�ˁ��l��#ݾ��E&q�.�U�����2D:��ԗ4�EN,�Ê��	��� �u��P8�j!�Q8�Q��) ��4E,O��NQ��n��[Ъ�!R� �|*��^q������ز θ�ԅX���(���s���'Dl���I�2�"�Q��e:zy��>.V�l~��s]ca㒳v{��٠]�$�=ڂ�̙:�%T���l�0����^��wH/]�\he�5��\Ij�����y�����d����m?1���.Z�^6Vz#U,��S��ߨ��5t�|3������myq�ZZ$\f̑��qf���K��r+ͦ����Ѽ	_2���}�����۝�,5G�2.�/AtqwF�t�R�\k�QY�����EHPI;D���IS�Y��u{w���}D�eCkN�])kyTz�[s"�E�J[J��&��j�_���E���i�+@T��;����0_�d*s�E�f�)>nr+��v=*����A
�VtK[T��v���pe7�}k$�.C}ʜe ��( ��/)��0{9����� 0^�d�z��&�>{�"#>�я8�=Pm|-��+f�t��M�ל*�Ǌ��N�'�=���&�V�0l�A����en0`pZ (o�r�K���������?ij��XPN-V�J-
0�4ٿG�v	�q���SQX�P��.��J�.HPpų0vpP����(4�/L�h����vu��.2N5p�uv����]�q�o�@ *1*~}����X�ru�n��ѭ<C��@Aa�o� Qw^�������/���[�Y��G_��X�[�[7�y��(��NS|OϺ辴�"$\�B�&�`5�m��/7w=\�4r��1��X.��?E�*��5�k�?zq
1B0����ӱ3���{~�邙?# P�!Z��J�x9)�$�������G�e�:����j+#Q�j<8����W��6����\K������CC��Q "�Sİۑ��B|�Ύ(�[��C�e�F^,\g,G}�B
���^.��-�9-������G��	ng�Z<u��ܭ�F�y�������� l |��܏��yGf�f;q��G�ctL$?$��%�������Q�^�%��Z�U�r �|�$8xL8����ƨ�S���ye�����(F�wJ�)Y]bP�C��0�(:�e�b�h����'�:�
��|�O��_G�FI_�֕�W�� 8��T��ۜ���}ۄx�s��͜���M�`v�;���E@y;W�ځ-Kb9�Ap�o(b�����aOL�y������3����_{�[���Ց E]���$��d<M4:/��"mj8b��|�l^�w2����j���մS�s#���pv�[0j���ń�}	����k�%���Ʃ����<u�i�?~�t(�� ;���| Cl���RRf��(c%�V�|ķ[�53���k�N� ��q�e/k�$6��N�d��s:d�]a2v Y���8_�8O���GO]X?�� �Oޟ���.0������~RCnnB��׭�Ɂl+������h��T��;R�xŏ�b펠H���;�&��,�eK�m��g�3�Lj�Kh Q�h;R3N�	��E�8|��El�IP�jh�'@��������9>b�<D�KbW;��Ky b��;��U�9�w���(����y�&o5W���<��e0_�,F�-�
������{�`�3=(D{�����:1�6��NP��\��r�����3pX{�T��u�o��g�+��I'&��ۜ�qZ���;��MV��Ԣ�Mx��uT�N�VSN���ԨB��.sV���\#�S�I�ҠhK��1,�B�Bg��V�Se��!u�Ľ��}v��u5Fl�gui#qA[��Cg����DNԔ������c�����oo��>}�՛۪�3�p��0����-z�J<`-�"�ݠ�ܿ���1��O�2�AO��t
Ũ���?"��acX�����u�׬�=ۧq��keh|���p���M�_�2	=AL,�q�b��2�Q̯X猶\;�u�jݿN��W92�^���@}T�%�K���6����&+=@1h��5�)\�Ӓ|CK����U%�ٶ���6�y�&���o�ϕlҲl+k�������߾���$A�j����t�Uu�J��LܮnK���'vDH�7<�	�Z� )Y�y!����O���F����e�ZQ:b}�/_�ZZ�_��Ȟ�SPZ{HH�j/�e�3��B�" ������gU]x���wջ���.��?�1�%�!��� V�E���W̦�~I�L$=H'��}�c�'�^��e/�ܙ���k�(��*��'��V��}�bBA�C�=G���o	G3]�V.���+�f�Uژ��8^UĊ"�����@�o�(�g
p������u��ZG�t٥���c?uA,�f��hgǙ�[P�?)������������=4������oFx��\�4ʂ�{oc Rc��.�;ڑZ���Z� �0[�4���X*֥���5;�;~�"�j��g�l�9�^R�4 �����q��3�v���s�Ζ��^�d:�'�Q���A-���)�Y5�j��s�/���I ��׎���4�`��gg\��X�xe��1'����A!-7�;��T[������?oz��@�.hg��[�����Ji@ɗ��x��D�
��p^��zʌ����ᥚ4K����4���럏���Z��Qѕ�(}3�\'�z����#o�Ot�U���� m�~2��#>d�b��$�L���+�-�F�~y�s�B���B�����3��҂Rlu�ޥ��'��>�5�	m�\�7
/
 7wՓa�E��_�R��ߗo�(<i�bU�ܡ�m�T�I���uNۓ&�Ŋ��l��o1�Շ}.�Pp~'�H���zz����b܂�(�zf
&h�K�j�!Ӣ�E�,3H��a�J�� �����5��g8���2C�=���&r�j�$J����̑.[��v�.�7222DGKO��5��{���DBTC�5���q�2{�h;Vi&�я�8ͱ4�~�*4��7\�n���f�@��Ց�ݿ���+��a9N�bu��WVW
����o��A�O��:B�a*���޽�aX��	]��UfK+��fS�2�:��Yq��'��"��O>@��~�p��<���R�*�/QZZb7<�k���-#�Ό��䖘�1��gAuufPT��F5���Fɶ�����V�[�����Q�j�n�׹�\�'ԝ��)��8�57��x��|c{�"�=�����kr_;��\1���PNB&�����:�t�w�Ȝ�	�UAJ��8b��=[��C������� vU�r2�ܿ;���D��P�3���<��*HE;ǎ�%&�f�c�h�w�X~���O&��-����c��v�jn� �l`�>xj'�+I��/�S�1��X��
�?�5F���}���U����c)|o�_�(�A����ZS>w�(o9�۠�]z���B���%@�Y�澠Nir��+�jF�}�G�1�R�鴂~�?��?�����4��#��嵰#��=���2���>���:�nHj�Sp�g?e��Ja��28,]E#_���y���tz|D���Y��/朊=��t���tR�4g����2��m����/w�W�R�>1v*h�h��&�k�����g�����^S��)P�f�ZHhsc,��ʖ͘�������	���F	���l'�66��eW �0A�ЗFZp�wb�T�����5��4�?\�-#��.���Ym���C��j���J�4������pZPT����0'�3~0�M�(�O�u��J>>Dr,�؀�]��[ �,�h G=���U��~��\G�E��^�\r�$N���T���C,�+�W�a޺��Ei1�W�K�&��g�Ǿ���#k_����k���+���Yvqѷ��Í�!�\w7�+��-�-h}��^���Ev8}�Ǻ�pfTѸt�x&�|�N��!���U��\x�cm��	>��垭�f�C�T'&.1�Rx4`8�3,�!QP(�Zf�"#Ɇ�[Zb�O `���g-���~���w�~S�A}�u���<�z#,��/ �����x�j�1�C����h�ܒL<��$�s�ݠoq�Z��e��~z�����xT���/�R7�da/e�g�5�\���$��1��o��V�;�E'�j�2̅IC���b��'�H�ZJ���
qt'���ͯ0D��^>��>c�M�n�����~.�%�9��\��B���Tm�U�h�t|����7y�h�Q\([*�ėg���&j�)g=��^���#j�Չ|�ڎ�EK��HB�4��;�{�Ebh�lyRj������ڛ����?,�*�\�AT�T4 Vnَ/Q�]��5R�#������o?{���0��jD>�����R��2��0��	��I�`���DKF9��1�D�N���k��$Ό�s6�oB߶�hW���2��((�*��$��mN�>��x��!j�W��YS��M�S�-ٲUdXy_��O��5ϦB�SFD�__�f�!ɫ~��,r�.�V�@����`;��(�8����({ N�nO��_�
<;�}�%\�gQ�}��J��?kډ"V���3L�(���PQ{�Q�P� ��K�:������bR3'a&���ߓ@���Tί��Zj��G�Tڃ������v��n}��k�?>s(��r�s��# ���@z��MH�I�d�Dꔌ̧;;k��u�7����d�����R6�j��}�U�O�׶[���{ETړ�^f�i�ث���>C���R}�M�^�g��!(T�*��{���^��������*Z��
���?�ۅx��i���|��+�۠b��$�9-�I�6 �7u��&z�m���e ���8��h����=O ��)cg��x`��.CB�2ڿPOm���?ў5����9�vrNo��W�-�^kr�>�����ؖ��-ݖ9{j̬����k��~X�3�nm&X����.__�O�7���+C�͛�5��<�.? ^�O�\e�O\<��%�:�߳�+�V�W�/|��%�9{�T]�IOO�ʜ��^�Wu�{�E��{�O�s�}���{?�@�E���s�ߨ'P�z��)"+��cBa1j� ���[7�JJ��H
~��yn��?�aD�B�~�%S�6��8�N~�?��ډ����r~��UO0[8$�g�G5\Ե�`s!�]%ך���.�H��κ3�HH]�^,2�n�ZU�AW\q@[�_Iۏy@��4w:�~^Svs\�L�.�-a���U-�8��wR�����1����ԚO����u����l�@�K��u��� �j�Y��쫁�NM8�ܳ:��u�ˈVA��l���s5����l�c?�т@��R+\�aȽ���)R`����A�`r?S����y��bą�ͦ,��ҫ�1�+r���ʔm��.+�� ��U�u�SG��p�J8��!Iv�����	s�g�O�u�cS��ol����*���@_�U�ۉ���e:�|��Ǆ􄷨�h������I�1���Ns�N�I�6E^U�Li�$�)X�9v)��Ȳ�oŌ��>����D��O<�[p�*/Zu��`?�%DN$���-�oLWq �)_cͩ����� x~��3oP���P����}��IZq�֥���h�����~qY�E��o�f'F5�o�v5y�979rlKv���]6i�`�b0�y��`��u�D�$�d.R5?̞�v�,���������n��'�c��AC�h��p��]M�pޞ`�5���̶�e���w�K���Ť����A�k}��@���E��N��c�ƭ�?�Ďl� ��A�0TJ��'�s/&�����C�jPv��'��Att6l���L˗���Z�И�qn��o���a�N�<h7.5UlƕI�.�Y\0���`��G��U�K/��9����K*�:�%.��R��-�[YoI�8>�Y�qǚ�?��;S\��us|��7'�oM���7
�\䁽NYo�찗E��^~�����w��MmS�R�,**%�v���c�hg�q���z����pW�;������2uУIQCrѣ�2q�2:T�?�]��v�Wdi˵�e&n�po�Uy�2�[0���uu���&�H���Z���ڷ�KÞ�ӡ���e�ٰ����I�kk�/���z��i��hk�49`�����A�����'��<�w�aw�;��t=�g�n6�+��,����G��[����u��l��d���ҧ�d6��!��������3꼍��>?��Ɣ@�j�NyN��r�I�p�Z�uK�)5^���>�:N*}f�ޔ+��jԠЧ���+�p������?�$��1J���l�aP�	����P�ד�a46j�&��� �1<s�REBx����Qt��D*�v�	�_���� *����rN�"�����t�����L��:��i܅����LwL�6���c�.�R'sZ�~�v�}�a�	��ޛ��+���d~�ȓ²������}$�v��V�%	��>OH�cf�|���o�@Y�?�9�{�i��6b��I��K�bw!�Â�Tz���86Q��Ds,�l�0�#����j3ԭ��p��'.MNE~�}ݝzu��O7M@��|�� �}T�M�.��Jt!���`�;,�!ț�O_�@��T<0�R/�P�/*���qϒd��~�c���?#J�6:���{p'_����m���tw0x+Ȟ��H�H��GvTC�t)pG��Y��c=�PN����EX΃_n3tU��q�B�JC���.��=�����eD�9�Gɔ>��T�F�D9L���|�ȡ���6.8�.L���,'��+�0?Л�m��"�G�폺�2��#�MDI�:N�f���i��oz'�|�B� �K�;y����F}2�Oo��}��X�X 0UCK$�����P�7��<��/>����G@�$5�7b����Ɖ�5�)�A�#O>O
74��y��E�M>Qw&��\��㬢�&g	����&O©h-���Ȼ[3��3�xF��	���d�S�͖���$�o�c��\6o$�LlX���^��&o1��?B�2��Zj*J��J�]�F�]h�j�����ש�I���u7��Dco�+�٫�Bo��Qw"�,X��R����æ�,K�h@@��-_cV"u�l�~?�s&�
����F��}��N$6_��c���E��ʍz��5E0�����ّQ���1j��-�&̭�G"�U��$�+#��w{J�?}=��o'�k{�c�+h��H���wV�C	��)�� �5'C����󳾸�&����kv��"K���/y4xΰF�C.F�G8���~����s.o�t�Q����<� ���x�)�f��6�@� ���QE�>h��@� t�����_z��I�L s�1�鸓��5IK�Mt�T�Q���� ocFz���]�i��䑶A �� D.�Y'C wQ�sg�\�J=3�T�$Wwe�t�"�7t���oڐ[A\����&K���++<#�Хs2)�r"h|ݡ�O��C����~[����ꮄR�A�p�PZ�P�\�'�r�:2�zw��<N����9P�S�֌�[ܿ_���D9}S�O�Ҏ+�[�X�6@���� �Y���WC�s�+�\�{':�W�N�e����2~�.��qz ZC6�A"�]�k��!���v$�5�7X��9� ;Ocg.ܲ��9��VC �}gp��B��{��ΐ��Z� |�=��oW}����?�V�拏u�e�W���� �p��bZK��hg�uR@����f��4���-�C���;Yb�~zE?!�R|������>!�0�-?(N���01������.�=��V��ƺ�R�<�E�偺�xx�T���#mm  )�Š���PE{���6�^��~�0��
������N����d�3���D�[X�!B�< ��߻9pՔe��X��N�M��������'�tW������[η(�)���=�|7�`j(�i4�-���cX�����.;	���O�ӫe���8�-%b7�͞_�$�vt�ּH_��5���Q]�����?�FP���9�e�m>%����Q�����h��1 �!x+�s"�����ط�?#i���L��r0��
~����H�s'�R���I]�g�N�5e��D�k��$ $/���Uw��M _5Ϙx�N�M�����\�fMK1GH���l�Y�����S���p����e_0c�����Z2RM�FR��򲃃���^ W9�u��/��n�8,R�q�q
s���E�Y;���oJ�:�t�a,��9���PL�Cm��5_Y�1�lx�u�r尽��1�)��6s#���'J�A�iU��u_���ꂍ|�����nyŦ��C�4 �ݿ���,���rQ������������#m6�G�F}I^}x�.8c�����*e��-�T �TM��si+P�!Xx:�	cn.�:L�ﮍ�'w��J7��+���c��v����%@"];�A��Y(ڭ��_q1U��l�(�NB��6��^cX�=dp6���L�N"��E�7U�4��*.��<i__�x�x����t2�~�"A���]�6�,�ל
"�������4d����]�0F~`d`�
�Y��Oİ�X4�_�W��M~�;;�}�o��-_�\�P^o����a�YșN��٘�����$E�&��S�7K��`J�W�=��}��O������$g��i^/OH�z {��A��ĵ�ʟ�?;jrM� wɕ��]OR@��t�4�Nl���֡���� �4��l�� &��QQ#z�W�6ܢm��h�?
�+�?��
4�B@&���N4~d��"�����r�r�MF��5G�X�'��M�[�h8	Sd� ��|��y2��`������4]g~C�;l'u�Lb��/vT�����'3�Úx���J�hF��J�U� 2q�S�3�<���L`�gHR�w�A��,>�:܎�.�t�������Z
����IO�H�]�g��F�j|q Ѵ&����@�����ߙ 'F��6`J͜ ��4��� �Q�H�1P�\rԠ;kb�;_Y��y�W��F�o?�h츜��T���Y�����ˣ@��f�<�5���11��Ps��`�΀��"�,!?�g)}2���X[���xpX�1�AL[�R��=��?@kQ��m�)�O��̶��O>F�'���k.a��ֿV�4��B���yJ�v���W��SF�"���K��*&n��P~�K$��]_2Nl���f�/-{�uE�8�ǥ��1��k�rAB%�mP`�DH ��'�y��y��?N3�E��{;�pv��	�_�� d��/�t��I����<�1��g�^��Q�+�2�b4�$r	��m�9c�[��b0yjȩe����14�A�	rXB��RU��E���:�Z$R��1�����G�۹�q �G"8
��#���B50�r(�C��0�E�TT<���$�j���fM��ɮ�y ��sR(�|�8��JA!�L-�	�9�(��K����I�b�T =�� y{'S����'�c����<��\��{?n�$�+HT�lNTM�I6��qV�5ۤKc�������<"�lLU�9���+�W�[!���t�@�Κ������$�@P�M�#?Qt~7y[����H��k�~��ޜrP�
��"]����������併��}������LoǣL���׶�JQ��)�[MF��cz��/Q�:��F�_Aw��{��wK� ǄO%G��!�'��,�ڨ���9A�c��3��1s���ihA����o��M�e]��7(��ˆ�h�[���䑡���"q��@��@B���^��N�]0��f��iҡ;�����?咶hّ�����5
)x4�YA���J|�_C�{�N�]%��rਗ਼�v�K��JO���C,Z)qNc���89�T�Q9/�����.�7�0*��'l��Vi���B�x�%��@�#�����z�qO6�-v��ʬ�<���y_ZS,w=��Z0��m�!=0����sG���'/Ɛ�E��Q��C�3�F�ssz'G;Hqs�s��2�y�U%�.Mv�PJK�d��ݭ�
���^kƮ�f6�&yD[�:1������s�㡒�յ��ŚM��T�Э�tAb��瘌G�����m�Uz�?�0�K���3s<�g���q�$�ֿ�3�n�Eoqԯ��5R��3�j!����Nn�]\rQ����Q��n��#�� �2\#�z�œ:��F����q���i��i�~�a'�*�&�@�	�c)+@Ĥ�Qݛܮopĕ� RC�P'�??�J8p�<��N���F1QL�tЁ4By����KI^�T��{�Jg���Yak��"���ۏo\Fߙ���^�����	.S�E���(����aEϱ�Jc.6a�_-��8~�ûT7���qa"��Գ!�cA�� "7F����k������ �$J-Nr���dҩ��-� 2/l�p���]��j�N#O���[)Q��q7��O��b7r���#��,;�����c��B��̧;r/K�5�h�Z���Ԓ9I���ef�1���|I�D�h��Ӳq�\�7�;s}8٤J�*dߚ݀�>�v�촭>�v�g 6/X�`]C���oL�{aT<gxiP?N�@m���;�72�<,�(b�6�-��(��r,a䝴�N}�$�g  �1P��T���R��`�Bl0L2���/ʏj�%�%��������޸����?w��=�x���e�ܟ�v�4E�aj��b�[3��Gܚ�#cu������>��|��h��N}���9���y�R��H��V��l-:Txc�*��M3�q-t~`	*-b��}mN2�ЕQ�l�"'��Z�����)��(�^m�_:x�}��åEE�r	�p�/����;���� �֮ߏkG �� �3	��e�G�{�_$p���=l�]��m�>Y_c��˪���`5$Qv�
绎�R5{_'W����w������5T�Y�����0��ⱞ{3B	v���d4!�;V��'#W`|��M��v,�R�zX�<p��6M�7w�|�m&sz5��1�q�h�LT�m��s'�\����w��K���D�:�n�F�v3#�4�+�@M�Z�ܚ/�j��{(=�j<����}�����{+=�������ӣ��sԱ�ML&�O!�Ov�sNи���h7�h_Z���4��F(�V�I�������:{�(2�Ip�~���%��ze�ԡuq��b����c��r�&���FFn���<�_x�c�3�o��b�ʕeZt�Ɖ��QAG���"��R'�D���uep!�)n��8���1@���kT���(��?�?4ЗH���t��=7�]�FJ�X�)3����k��򞓄l����U�u���~|"�=�[Բ*�6,\����W.N�Q/�\�11��� P��{BXZ*=qS�z+������,�
��ZP�v����z�^�7���b�.�����8�R,���I��o�d=,�A_[}�m��>tpȶt����ɜ���)���/��s��<ٽVӈ��i<'���ViN9���#�rx����<���]����B��(�ҩ�KM�
�����_zh��h��/�@:7P��o�с�e����4�M��i��ā}��H�m��q�so'۷���P�Q�&'�!�Q09��N��G��#u�
����:��\���������C-��ޘ#�c܀ț���z<7 q!�1��Ҝi8��i��f<ƛ�l�I�$v\�m`�3y�Τv��V?P�'>˖�{����y�+��%�1�!^%AZ`��pIE���}�^'H�1������7�I��X�&�%�SS��v[ +�F���B^q��%��7�v�!wjq=k�봓��+|~��+1�����힒J{Xg-9u��8�$l�zk)���F��
���W�]�"�*��+*Xu'��Q+m�`�=q�E�5G(��p�g��9�gK�b'X�������3 ���b��O��.�{���V� {�Έ�C��Q��;��˔�Q
�H��:��@s��Ԉ"|�#�C0����PV)�"���M�N�Ej�E��u����!v�a9*�m3�|�s'g�1��p�U;�@���SB����o�<w����[���(���c�	�cnPw&<���~�� "M��� :�'��|�ה��"u'�NploN{*�z����J6�jw�A��n�)�4�S��4,�9���ɣ<���cNo��&�����!֡�����t�jC�6��^�cc�#l�{Hw��Go~�����q����8}(�F�gW�y����{wj1C|�(�A�B���^�~�+,F����>�!�	}�҃�=͘c�T�Hg�v��a��i�x;c��H�-)rݑq�{&�?%��Yh	�܎�Å,kX|f�&�ϭ���s.�A�R�Î�Ņ�N x�Y�'�u��,�mk�We��L~A������?�\_�z{\/�&D%xc�˸����/���� e?L'B�����4W\g'��$��1�n8>?cյu,!�E��G4�KZ�E�b��:�v�*���Y1�P�&�9.N��P�Yc@�-ЉL��w�(%n�E�Cz;5g%o���Tv]���݁��\j�	7�����HUٙN+��_��ٚ
 �+]7(>2��% M2Twz�V��N�pz�Q�c�.i1/_�y2��A��^[�u�ih1¸���,Y{5��$�|���%Wޗ!� =h�;��m�y��l����(W�՛7~2�/r�/�����l�~<� 2Q@an>EF`��@G��x��lo@:p?'%�����p�<Y7�A	���R��R<~��%Ÿe�="��;j�HA�V.oC�Y�*�"^Qr;,�&e�xY�|�bW�@4�2.� �n��ˉ�>j���z}S�WZ�c?�?j+��zS�:T�ъ&u��%�O�]1ۏ��#�nZ�Ϊܧ�D��6v��g-B揫�@��*8�6}X&	Di�kD ���3��u(���9����Q��u��F�C���7�5G��G�o<�k��8�����o'W��#'�.�m$e��1*�<WF����� �9���	�|��3��)1��Ձ/��x�ۡ�eI�dwX`bO.������$^]e�Ũ�3�[�������'�+Iwh�m��7����m���F$�؍<��w�J�l\��P 9�̣��%���1{Y1����Z��usI��ќ{�����gV�4sOMM�`��IÆw���(��3��΍&���\2%(������V�kZ/O�Ȭ?��9[ѻ �ۇ�+���y"4r�r�j��xl�6�����0��ņ��>aw��I,�Ԙ��ͤ���� ��k� �t�tI
��R� �� �K��!���R��%� �t7�t�����~�ץ��z�<3w̙����+�/�G�}�_�z��u���ߎA��]�-��J���ǖ�G�l�og�ד3{�ǏՓ�J�E�l����R��>�����x3W�ۺ���}F�hc��.#n$�p�^�[�&��}�9u�r3�H�4�5=�<b�s���I�W�s�N<�̠X�d��l�˔%�y�.�7�1�e�XWg׬��z�X2�X���ڭPQ�����I7u�5���W�+�?"f�~)c��'�|a�g�)&�lH=5'�	���ȟ9 ��a0=���r>��nx�觺F����r���<l�Vt�LS�l�\�Eߏ�������s�)b�bXL/.ל���碩������X��mq�Y�H�x���e<-�����������zV��zA�R8q��p�m\x8��oLL��+`�'omXU��L�!W"��w[�ͭ�R[Q/?;�<�=�
F�ό�d��*/�Ӝ��A�\���D��``�u�(����,y��%w��Q��u�?7:C8��ZIRp��	���FFD�|����r����7�����ވ� �����P���w��9sq���O�h��sG��e��V�!�R�%�#�P.o�t�_Niu��w��G�'�@E�C)���?��tu�LX�o���u�l&'x�HVj�C|eE�7�)�|��0�����H�w]2޴i�SDNm5�C��yB��/� �\?f��"���Tz$�"���Rgʹ�L������vC�ֿ��v�D��=;X�����c�%p.�g\lj�x�Z�g����b�#�I�R�)߇�V@|���L�MO�Pښ�S��h�H��s��u|�)q ۦ�k��Mؿ����|_�J�0���m�C��~�%�
8�f�;%|k["�	߮J܌Z\�𫃎������@��&�~��0#�����S ���kwg؛r8C���Ԯ�J���F��g6�%°�K���KϛZ!C�T�0��hf��Z��j|���O�V7C�w52@�\����{� �0���W���S�P��g�;�=�Ѷd:[���d�K��6hE8X���,��ܹQ	a<���>5���R�Ss��x� ̍ �빑Z>rBv4��q��߬���)�z~)���� �a���h9j���zش9��w�A>!}�����3 v�����Q��' �	U�����r�9Xa��P6u�y0�G��7U�����a��Ӈ3]d�������î�أa<޵2�\�QW�x(�sj�=pAOGIv�),�����a�~Q��i��a���I�=C+�ɕH��3��`�'��ޅ*��=��v�7�甼���7�/)���s/�(�S��-�$x����^M�����+o���ʊ�����S��TDo�r��)�☚��TݽpZ+���f�E�L,<�.��2 ��7ң�j���D:�q,�:b���#��|S�/x�M�v7��`;��-���gcւҮ�b	?�!g���@�/!���5J�в6|p��mט+%9�O��>�Y��=�嶎|� ��}o��˒����5Y�l�t�5�*;Gy�_��w[�8�p%��/��CW��Z ��}U��ҿ�B傴���ځx����D�)٤�n����Oт��A��nPo7X�缨����e[����.���Ļ2�4+RI���"��è�Dsޫ��2:˲���u���Q2(g>�H!�f�yu�s���������<DnăKG�³5���QCq����O��bQ5�L�i"�������3�U��o� k%�P8'ɫ�����'��E�!�<�!��Ѫ ԶKR�{s���O积���/XNmg"���VA��=��s�8�1�.B�$b�.Q��29%�{��G����5f���n7����%�k��.+��}�}�`�����9}���k6��K�jH�2 Jb�X����	BF� "�� ������q��b��L*�>Dy��/��k��?�Sz$cq���E5I��m/�s�	�3�](g�֔ֆ�P�73�N;�m'f�3Ԍ��y<b���{�����A�?�F�-1�(���%J��;�%���j���\'WR��=$�;�AIz,�f���a>4x����̤�e�c�2��ynT�����$�GF�5'"e�'o|�d������'~񔳄!��O��=���.�f:�Clz���U��Ywm�Pl�v*�� \�N�ҥԘ^yu�m'�F�Y` V}�����U�#Y�:~�lI}�к������#�#��:N���$n��Xh��;/�kjY8d��w<�~c�����o_�ts>�>��Λw�9)xDS��я�P�
�W�A���Є�p�"�I����V�CD�H$�����X�Z���z�lc�3?&H�����s�],>W	^��{��|\���DRO�98Rn�xW���2Ѳ��@�t߶g�U4/?V� ʐ|m'��b�A��gy�nĈU#�
gr\�v#�nt�<|�z8�ƛ��$��NS�F�����;�0�
8�᧯�Ya��h�GP+L���@�N��\="| h�[`��P�����E��鸆L��t���l�7�	[JW� xT���ir�\w�,��^��T|`���"�N��%�7�����ݒ�����]f��C-�B9�t�7䊗�t��L�S�V^*m������������.�ۡ+p���x�uC��2�jZ�|�ڞd��w{�"�Vڸ�S�]?�������&ܝ�5f���n���-`�s!˲���|��o�uf3��I�T��&x��'H8/O�d��8{̊��P��φ���'��u*R�k��D���9#��.� 	����g"R_�^��)��>p��(Z�'�j!���9�r�=kvq1�����$i�O�V�7+~��M�H�X�l���WV��O��}yY���ۘF#�<9�)�跾< �`l6Pֈ��)��.;Ji�'$��PY��0@�e|B�P{ϓ6z���P��`$�f��p�����*���������C�\r�wdb9X{c�R$��]�|�SpH�P�w���a�c�h*�#F��z?�,��U�%�8�2�,���Z�/F�v��W�!�$��O���-3����ۧ��p�#xSh�*#����w@�1�$E�K2�**��|�FF��1��5�nJ�lM����rFCi}8�B��!��*P�w4�I�k����U�`�yad6���B!sq ����b�������˨B��=���f��	v�+_i�G��j�I�&�e��0O�����l[��Y�١:�Q!�~�����Қ��#1Ԇ#*34�r�,��5�����`X)������3?�WJ����d$�@5��<�R�(��KO1]�}�gh�
C����V��䷽~��-���ʆ�)�4,A�d��4,ϻ�f'�����Ջ
�R���ȲL�!�����>�#Md}7�hd�X����D%�^�D_��{:�xR�p��Q��4��*�v��hxK!�tEg�#?����!�>��w�ʆz�K����8�F�����&}��B��}������ٝ@�y}{���˷�C�iO���Ҿ��>|i��ǃ�Ԗ�6���ެ��c���!9�ǥRt��p�ecaG��T�{��p" ?6##*���Z�硚r{�ގ�=wJ/O4A,�9�欫GT���}ĭaǃ�m9�<�O��*����A�-�lI��ȴ������ <n�xH�|̡�J�ПY���zD����������t���pdcʵ!�I�&���Q3Y��bg�^���@��F\�#]����g�P�+(*|(Qj�x;���p���"�+� ${�l��;��E;�§�9�-'m��Q�j�Ñ횁ǖ�^X���'*.�Ü8��u�n	��D?|_�<���K1���v��̓b�g��b����p�����w"�l��Q��T@����=���;(�E������(�Z��;��|���[�O���E޳N��70���n�b?QI�[���]֭Gq͇4�w@��a��UՠܯY�PףM�ć��+�.ǯ$:������R� � ���vP  ݂ �L��Z����(�[� ���{�Lb��<U���\�����ȟ����l�̍/�,N��02&�:d����z�]��C���(}�C�իbU�<�|���4]s�}����Vk;�]��#��
p�P
jA�{��aGě�=6b(�Z�в�����?j��l���"I4@�����> n	f�><��isIp�V�*�?�WЂb�����S|"J����)�j�n�j�2������G�g��UC���`�������z鿡��|o�(��u��Y�
 ^��C��!�J�� ����"-�d�����-eۗc���H$K6rƿL�'��q叓�M9��/��((��+�ؑ�P����-�K��Q�l�_:�#��_�X ~����M���^ʐ�΁�E�y�K��5���R�k�T9��fE��1��� "��C �0�W&���/�g���Ն�i��C�Ym��2 ;��4��se�����#��|�m� ������ľ�D�{���l��������Py[.�?-��c�G�G��֘��?��Qc����2'Wo��x��ܲZ������Sq Ֆ���y���H~����"N�P��2���`�Y�p�Igh��3FQ��u��pv��E�#���R�4��Tm��dA���}֭����F�k\Jw�s�J�}�c���=s��8!-\#	���s�ԉ����?��4@ �C�v<�n#�2�ɑ��wT>���7�cr\[B45#>���,ԪD*���**�e(�����e!�>�l���>cC�}l���q�Uß��m+���?��Kpr<P��X�Lj��B��L�2�J�n�x~�_8a-�x�37�L#�4۳= 6P�_�#y���w���/?4�	)q?PzS���>
RT�g�i������c��'I/౰�j_�^��~�Ė�CZ��+���C����-���b[�s!\�F�̸�b����r�K��⑭`�ѻ�<��D5˃a���4�P�˨��u���7�[؝�r��`��#�]DM���ȁ�8#�`��s2m&��-�4\s��:��=�Ž�W��j=���.��9 j��멹��g���������N� �ՠ�4��K�]��.�vT��^�\f����/ܐawh4Ƥ5P�)��8�j����:�t�կ�>	�?�c,)���,&�%<Rx�.��X��[
BV����/�p_'�

�8������I
+	il��2��9,�N�}��1ȱjRҜ��e���n�Tt.��<���t�v!���=���ߑC�^"�!҄?A77~L�$����)����3��Ѯ��'r���y�`�x-�vy�z\����栾�������@��/�܆�1m&�r�|��Ы�i��4pA�e�)V��!r��% 8)���qƂI~�zX
K��̋����
p��#n�_�U�~6X%�'���
�5�I�٪0�v�R��O]�U��ۄ� ���)̓����T���~�w*����0	�$�����2��=%���8�i����/
�XH@����,���!�FNy���N�M��R�D�߉a��\���͑u� �5�̑z|_Im�Y�X�Ź���)�K�p������A7�}9
�Q�|���W�����B)<p�Д�4��c	?��<}Ӈb��l��h�~o
I�V�]��-(�J�N�|be�g�ǐ.{�JbS��t������\��(_[�U���{��E��_��i��ǈ��\�	]ܑ��k{�"�8_�E��Z��N[g	�ew�!]\D���$+7z�so�Do�����⠹5QMgJ��ꆑ��\I�?U��πE��)��rY���r3ۙ�FSJ����洼&�	�Wd�Gx���@�}�\Տx[쐣I�p�uj�2k��c!	I|x������	r�ی��Ƅ�G�����#F�0�Y���+E!^dr��iXU��gG�9@�o\1� ����S�o�Af�����-�� Q+��e��En ��vR4p�cȟ�1�,�b��s�{~����r���/R�d ��բ���/�Lg��6o��aJ�1�\rvƯ�>Q]8v|�f�Q�xIT��f�!qy�T�D�#���i�s�Kߜh�&������$��G�1+I�cD�Ib#t\��v����% �I�~�E��;>(�l���������N~��?�*�5p�&Z�t�>'��i�Z ����{�9ldKz6c;�`+ċ<��� ]q��}�m��WV3���X�q�
#j%�߾���s���=J�8ɫ0�>
%�A:��U�]��k�Y��U�+~�j�I���~T�*����1R8,:�|\�>�]�?i|Ɨ��̲��l�g�}c�!�R7�����6GT�Q��V�Y$��B�;S�ۑ37����l�c:Ŏ��p6�u9�f�8��R�{�>{�4��&F��˄ܜ�U^:B���3)e�V�0�3��I"�;iU�:T�B�]z���$�mԄU����E?ɂ*Osl#��h�늣��@��z�KB�}'��ȵ쮃i�'Òl�9X��RLwf�y��|u��,����g�i��Hݸo1Sȧ����A;���]{x�'�
�C������7"�$T�y���1E�u��9��RV�jhޥ"�j��y�y�t�jQ��W_��f<��u7���7q�ȝ������#C:�T &V���'���l|є�s���j�{!߾�o����g��,�P�I���/���G��i�9u�"kӆ� �˕U�$g�2P���J���5�,D���|.����u����uq�C�����c��y��N�ށoX��+1KIb
ޏifj_3��#[���c���/��^|�>o�p^̵�e��u��t`o�#V=�D�].
���gg���q.��P�e[�Y�I'�N�1�!``�A2����Q�~$ZNQv�~֞tch���g���ۥX�����c�w�6�m $�dqBZ�����h3D��޽��_X��D�7�Z��Y�_����ɂ��cq������l�D�S؆�̠Β���0q߶�0j|�؁��$�Á��\(��O �ſ�E��D)�5�}ڌ1n4���ʠd[Mi4t=�!^H���b�%�hV���N��G�^� �-�M�~�ZR}�ء�E�|�Xh���!�wm��z{H�����C6�,i�j�a�!Y�-��=������,:��7�jhəv��ʱ|�l��K£o�-X"�mD�s�	�\P�S���F��m��?3�
"t��,��Iǘ��̾p�����&@~��ZD�0���]L��M��=���l��Y����P�"��AD�+���T8Z6��� R��u,�r>3����w؆�������26}h)�g�pHd��z}2��+�R*��p�Ȗ2Σ��1@$B�mBO!�&�rɻ�r�K�աҾ�����~��YȌ��>�C�o������2B��7�Ή��	R�<��pz�>�:5y%�$|G�4����*�;��`���!)���S(f?���P��m�)�s_i^��:��2�#Y7��D�}9G��|n����&b)���G[}.<�ġx}G��|�g���������j(�-��Yqڮ#蓬W����^^�LY�N.��ʆv��
�l\�B�&z<�G�Ds�Ԧ� 9�/�N�'�Gn�#���Y��JI�W.��a����z�l;R����Χ���@۰.m.l�Dn�u�3$r���O4V��VG?���ӈ,�[�gU\�8��^W�������p�d�|^��4D����Z���
�1��t�J��q�Y��7Јbb;��U}��z��!�Z���}t��h�\�x(���,~�q�<R�٪z^J�M�(���uu5�y���.X\p�˹Δ�z/��H����X8��k���x{�� �+�����{D�u�c��4���w���S�M���+��t�����G�}�Y���YY��茔zF�ҝi.�a/��U2�Ly�IZ���t�O���Ò�d��˔�Ƿ귏�"�e�=�±#�X��i�TM�s��&�M!�.��{���Bh�ɩAJ���b�W�#��r7.`Ʒ���ڀɫqBV6u4�$.9���~�C��E���;��J����<�*��;*���=�u��R��a)��x���-��|��( ����wJ���#�,&�BS���M k�d�|�2p{i/��=So�#�]ߖL�4�Ǡ/��}�{�8�x![Xa�wz�
vz.l�=��YjV�Ռ�?���E��8x~�!_!̅��p������U�C(/�{dY]����NV��H���P�oZ�eO�ӱe
7>�#���� �E㴜P/��ϓ�u�Jn�tM���u���S�?����=�n�LecM ���Q��>��ld��&��̈́}�=�Q���*��C����c�tE�0�,P���U玌?Z�����'�1�1p�^��JZ�W��e���M��4�TGxU�c��K&_�Z�L��0������)@x����
�E�-��3��r4�+���4ZA5�
,�տΈC�\
�����}b�{�b���w�(��Y�v�岺��Є㾳�Hy�R��#����i����"�S�3��c��M ������3����
��A�,�Q>S�5St���~�
T���_<����w�~�+�NзR�|�y�Y�<�j˧�K�����4i�Z�mqƣ�tAW .��^��p��z̅>�h���<L�Q�)Y������C�ݱ�ki��JG�a+6(T)�>���;��G�|�Lmֿ���!�YT��s\���ѳ|�e�O�\�UU�+���1&������S�#])��������K/����.c$r%��jօ^�]��d�-�S17��i��vf��Fv'ZP��<qj������/U��\jB��-vN�0G�
�&D�xD7;(���êp�x#�puR8M�0[ZV_�seQ�M�}�"���͏R@�M �i���Z�l������־՛Z��m�[(3�o���Od��J6!)Gg�ۇ�|����T$��;+��N�7��=cF��ФƸ-�,�6�H�d#:��q�3=���,����ݞ���VY����P��g뺉�1ZG>@� vP���9�"��b�J��솓	ŁrL�o��!�ܞ��k��e�#־ۚ�ʀV�Ջ�nˌLJ�v��i� $�w�U��Y�Q����d��lb�<�e��/ih!ĸ(�UP��}�j�Hx����`��#�*OMg����(��{B��=e|���!��F'�n�h��X�^X�L~a�%����8T�&5�<�:RQ'm-�|���,�^$�}��x�.J@񖥩G/�/��'�Q�E�2�%u3�QH�ꀤ�H@I���ض��C�V�eѿ	d2��_Aj���x5�P�sc�ݙ����O�\�B������'����\��?^�=Ѯ�����/1�����j��(��m�clZbˤX|SZ����e?<����ʆ����km���Z�I����@I���כ�#6<�U'��%��U���M�$P��3�����C�Zzx��HG�GXA�mK�d��9��t�h�c �Q����lt�U��8E�=�q�����J
������ ��h_7�&K�ks.����ר��w�@��J��(�h�.���lVX�C,����R�pe���$n��3y�Kđ�'�l�VYp�bT���"�h
3\�"�\��B�HƜXv���vB�Xn�+-�֑ncI��Ф�#�o]�Ur2�n���[��^#]�l殜�m�wa��ůJ�3A�f�q.Y�	����[��:�R�~.�_)>o0˶o��U�eS�X͑;�F������k�8���hA�g��k�m%�T��(i�(�z\��r-��^Ǒ�a�6��VN���߾��?q��v-a�C+^>�@�AjPHK���)T�8�3B�G��C���T	�c��"��mw�����F����[|�≳*�o��u��P��oy��@�A)iܺD���݊mk�7�S=2�d�rE�B�����k_Q�� j2����LtR����"������~G��X��V4"D�e;�y����4��4��K�Z�E����X���CÌ��1��v���_!�N�3�֚�"G��*��'���s&�F�jaI��F�O~臬�B��-���)/-�ۈ�B
� �J%��P��z�\�7X�^�Վ׼�_��N=�/�7!v
Qc�^����|'�}�<�յx�S7:A-���,Gr*U#�W��-����:��cw;���F�XK� ��H�ȩ��m[�K+N�q���}�#�C��27����6��͌R����?��7�TMV���4 ��a�9���kc�r�z�L�0�aT{ν��8�UY��e���8PH8�1P(��d`�iyM@�+��5r1��&�&�ݯp��"}q?R��� Ӊ��8�ƿ#a�\?⠣�*&4��	�2� �JG�r��j����;���I���>��ֲ�Z�X�
����I�t�~��n�
�Xb'�I`jH��[=�8��tCTɣU�Y�'��pp�wj&�s#�o)��y�Ó��p�#Ȝ�'+O���(]ޢKl�!0�"�d~	=|oe�R�75���p��i'?�������őh	A�j!�E��������2r����-���5q��/衫�3q��F�-K��`���6����eL�6�dafp�� ���da<�/�٫�s��Z�(Q�
%���Y�ɚAg4���hV=��%��6������sӹ,t�^��g�]�����;��R\�a�+,p^�����IA����Tß�Y.��8.�OJB��GJ<?��&HZ�5D `�=��&Y����N�G�N�F��h��;!8}�u�<+����3�Hb�-���p�n�7�rK�k>]�=Ω+Q����$�,�}�͞��j�2ॕK;b�#�MR���S��Ֆ�j-:�r�J�+��l; ;w�L/���������4�1��y�X;�1��T^� �����2$)�(ڶ�D��ma �j��:���^�^//��lI���~�19��04�����8C����{��[1j��"B��r����V�z�	�V�����C�=�����5��}��$j�j��!G*�J:��#�aۉ}���~��/�q���Z��P[�9��df�۔���%�(�&z����o�� ;�C*+�&g\�(i_�a�Դ)U���<4��J)����� C��8���q�p�YPcŚWɄq�:��R��n7�	{�K=YDw�ͨ��>��J7cu�_3��Sk�����y�3l��۴�f�1�r(}HܺL%
��0�:������$Ьt���YHF��lM���;�K����M��8���6��`��ON�o����~w%�+we={x�)џ���a
�<ip%�+U�dv����a��2.j��l��8b̐�z*Qw�E�D���!��_~�!�L����x���'���PG�����o�T���c��W��z[>B|�\����,g�1X�R��ߪ@?�9_���v�K����8X쮎*�+	�ڢ2l���s,��S����� <���)q�����Il��!kR�1B�]m��A5��豽�߉�G� �Bt�d��QN�Z�=��n}���8��I��6f.�����z'6�RM˔��@�!E@�4���>c�XX�C�Z��M!����q�uu
���l��&���HՁ�̈́��S�b%>F��Dҫ��)�[Y��0*�W`�_X� �4����\�7Z�C�G�m����;���|��;l�Eǰ�,� \�\_g�9�0O�V���������	4Ķq:`t<�����t/[���n���0�S	�) �H8+W����M��@�l����-87�Cl��,�|>x�e��:����h�C��ٸI��8�o���Sr�/O72�N ��%Z��Y�UM�Y�;�"=S��A��ąz0)�|~ZA�?=��e	�act���n7���;�8�󙟃ru����#�D %��?ꧪ�g����y;�¾�as�o4��)QزB�ps�I�au�VR�MC�7�]t�W���`������G��Sϰ��$Z�To��+v�:��e��&�C�q>D���p�U켂�	�ȣ�oG̟��Т%�}�L\�o``�C���vo:��>q����\����d��=1����U��o�ly����z�2��t�+�7��%Zrw/�|��ᠠH�{�Zަ!�'��IR�J��x�y�x)�P��J����"M�j�"c�@�b�����W���`�#-w�K�r�;�=��Ͽ0 9"�@GWh�;�9����U؛4��+6�?5c�WG~�<�Ռ�'���M�
�o�-�O}��l}���eFAb���"�I!#��_=��w7�ߕ_e�J���&#R-ȯ����d�P�xi���E��=ɕ�#	n���i�l�Q�BW���~?�Η9Z0�y>�{��v���󺜞������K�Xp��J"��C�@�����&@t]6��#	̊i�X�yC�48E����݄��h�n����?o(�,���]O���׼I��xCz���/�����׿�O~ �Q�Jޒ:k�i�<�D���L�|�P2���RW��v��țkC'��3�s�*}o*�~~���K�[g��y<�}X��;!���ŭ����n��3�>$�t����S�Bq�F��4Q*��X�U�od���@����W��Aċ>��(y����[b`���)�9�b���
[�V�J�
�]M"�:ET��Y���5�$ѻdr��Q���(��#�� ���5��@0��U�jIMV��E�:�E��Ws�	0	i�Ǿ��� ���S���L. �ib���h��?<d�P�
�?�y������x�;���_�+�:@]���������θz�2>�a��G���c��o�`k$�O�����);.��\�B��_؛�b��#8>e�ی����L~�^IoJ���4�0�>�RϠ���"�}�Rn/j��T������X�����D���1�^b��I�k�!�Ǖ�������*?;�*9�$	~���֜əUG�ڙ�O׆��Q��d�Q'� >�Pґ*=V�c�I2���}���HQ��*��Ux�3F5N/|�"��(��nc�ٚL'�8�����o�u��H�,c�����1�7C�D��3]�>|[�=�)�Z����"�[�vh���Ԍ͠l�T��$����\��.}�2L);�7K`u+Oz�K^H~�Gv�S(��1��ϧ��9<Z$� �2�^jn���i��p�ɩ�^�o�� ����	F�����u��؛ĵ���OZ�5�$O��&)��Y{�E=b���$9)[]�0�S*$��o���޼{��%~}E��5PR ��#{5m*�S���n ܼI畦���g$H|#�a��\0���/��_�D|S>p.7m��ᔤ 4�'[�8�Y����3��U��v�D/ɼ��cq��;�"���-�E}=.��F����ng�4�8�I@)�gh�=�r*;({�)ə~y�f��dhv��������ԋ�=�Lw�?��9uTy�>0����4zQ��1��P��*1W|�a���d[��{.+=�Ip�=zGׯ?^m�'���q�T�c�	�l��X)k�,k~e��l�l�H[�l�bc��t]��h��9�h!F)T���ە͔�Ǜm�6ƿ�"�T"��F�Q<�x��6|��U����Q^e�J��6�b��XMs�z����/_�z��=��*�I���X����=.����@F�P��J��=��YQQ4�OU"CS�t�S[��k�TG������E� ^�e�VBZ�LTϻ��+���͚+���Ë����DD�j���� Q�����K���
�5	K��Qְ�I��������o!�~X��Ԁ�14�'0���2�~�r%�7x��`c��Ȭ+�����\�K���L�<�����J��Q��p��(�k�J_J˗h�4����h�p���#䅬zX��V�㹱uS�s��mU���c1�YY�n#����yS����������*G�w��5���ݗаj\�H2�{�N��+��R�ya�J�r�q*X�	#�l�M��j}�a�d�U��S��[�w�*��Y	����oCDh���zoyU&�b1/����l�!�9�Ǹ�4g��)��f3�������OO5��+x�[�% �=�ѸbR)�֙w����S%/ƃ�څ8�xU�����_%P�|I5��g��?�|�W�⹭�;�k���$BN�O@�;��(q�����D�o��~�QzM�_�-�)��24t��]�`��m�_�흎5�V�Kg�J���2�Ci�xn\n�f�G�2��ʇ�D��_�F���J_�:fU�qm�f�2G��FeO������DHu���\*|f��g�ݻgt�Y=<�h���K���"�U�4<�ܮȽ��5Y
QJ����+k���1�ybh�9��qxe3W���Tr/?���J�x�[�␺i�MEm���j&E��`X�/l��S�Ä��;�V�1�����Ξн'�{��+?�j6���:�_��c�5�7����9Uʁ{���s9����T��Aƺ
>c'���jT��e�RCƦ����Y!Y��p���?7l��?��DI�����\���Z'���-�I�>�I�UnR�7\��5g�����d�=�sZj�R�7�W�#{�@�lׅ�p:�7�e�7��j�S��*v� ��F������y(�Dōz�gesɩ�����Q##$�n�钴TO�Ms�2li��>I+�9{�ED��~�-g�$S2�OS̤�
䍉��d��e�?�Z�A����	���}.g�2������X������o��s���U<k�8�'�q.������&~bv��ўc�'E��|��^b,<��0�ՠ�ޕ�׼ �2�!�#�4�v���3Hn��:.���^�p�h�(Z���ܷ��%`Kl�Z�s�O	���~�z�Z�M׎�p������S9� ZY�U���J>�C.�#zb$|	9��5��R?�l�
���]��	/�ٟ���`I6��^��r��<����mX@����B*4	��fQ��hs�C�D�f��Ww߾����Gg)i�au�<sr��*�;1���#�&$�
�6����?�������+�j�XIM5�x��<B^�CJa?[d[��ںF����^�-K��J�4�l�S����k�P�\�[��R����#�.&ƳV�Oú���Ui,�(Μ	���,f�#��ʀA	@�������;,5��CrAq�%�^����JWU��6�]��/}K�s���^��C��}�V�N�nI��k���f�d�X{�&>���_� 0�4��mX�Uϗ�~�J��nYĻ~���O��л���w�*4�e9�>g	4�?��H$��ym湧0v^�f���&-P�LY�\�췱�����&U�x�,��EJ�N�P������|����/39�
J��������s�x�q�C��hm:(���A��Sw���BuQ�y�D�LwL�O���UE*��}[�ż�E�p���b�V�G��m.�X3pܫ>�y>�%/Á$C�������W&S�����/ԝw���0]O������D�o_f:Ŏ��P�=^P����Q��o�Ȯ�Ѵ)rkkX��^�4 @� �F'j�>Wz�9h�����߶�該Q�캬�I[�=!�l�����_�ƮM8j�xL��Jՠ+_3���r�ܹ��-K�Y:q��(H����r��2�j���5?+�%G>��� d8��qI����-����"k�g���}C R�`�z����oƮ��_®�� j�[��w�+j|�n�@�d�Q��pLF��g�4DG�߶��犚��+�Q$jn��ؼ�,yMt��FX���N�jz�o#�H� e��ٶ����[V٧T$�ܱ+lU��?��A� �����ߎo?9���g�}!v�c\z�i���qq=��&�n�F����y�&]�v'�H�:�1-��Pi�9%�
�o���,֨(r�s�V+��{�~Js���/1�=U>�E�W��&?�9R�&|I�V�/֬��R� ;�/�hEYʋJ�~������j(b�*F�C�uKRk�b�/��s�qn������w׸P���d*<O�1m�_�$���b�
D����$���(
�����ˆ%��8��_���J�y���U=��+F��x5D�V���wi�?k�R)�Zq��y���������-ZNZ0����ܬ�h~AJ �'._b�;9�7��p�Mo�y	��#�rtū��:6������	�S�j�._�~�MkGP^��w������uEd�r(*0�B���)^L�BVP9�0��i��=�uz��)~�v�f�ZJy�`��L��}������!]t��U��5�	LR�o�Rh0�((��V����wF�?$<�2K w|�5��x��:$P�dZ��{1�0�im�dR�M�����p�0�1 7��WJK��o��*	i���j ]�k9}��}q�ֱf���M������%,յ�u�Z/������N�a�[��
��HŢ�3=�x��6�:�o�E&&I�����j�}���UϘK^v��kG��hn��m�Ӓ�h�X�8�;Q����߃/NEW7��)��i:��C�y�|���$Eq�L�WaOm�4jYT,� ���_����BX��Ң�[���`����<?(T�!��vOcĺ&��n$?���ְ~���PC�)ďE�?{$�~�KS^���_�=)�"��� ����������^����h�d��*kZ,b�s@bӃj���:(�����[�?C��܈�C�A�����v�:i8�3�@��!?{��︅�챻�1ä�x��_�&lK#���W_���=����������R2�R�ݩH7��R�C��HI����ЍH�t�����f-��0����O����7o�'{DJG뻰Ф�`xVVYȮ�?�	��W�����k��H��ϑ����k��N�(�;�a-6�H� ݜ��TT�Q9`xIdӊ�I`�RшH���@@(�N\�w�LK���:&�T�L�&�c�S��0���z	��<����[U)}�w����<U�y��Z�L�t���<lܛ��|h{J(�k]lp�}��V�;M��*�'@�e����ڀ�gM�gF�Ly�j!>I>�����V�����2�U`��r��e	�~�:�TX�{�U~W�`�հ�Z=4Ht�h%���*g��Ap����鄝�O{�}\�A^Pt�+"�凵*�f�v%�HW����j�y�� ��������K�y/%��ޅ�پ~8���fO���&��É�M��D�B0��k��h��qf�I^n����[����'�
�ж?y���5Uwx��������y[�H9|��Zwjp��H�]�����(Î���׫�i/�U.	��[��С�`U��y[ۖ7)hGn͝�Ue��S={2�)���K{���F�?r[W�����2�����YK���<V��x�>6\Iot�Mq9�yN]���ܰeB�/��$��Gp虄���0����+����4"[.8�*�V`�Z�B���Ք�е.a���|�)�a,)��:6Ф����]��C�w��e�OP�� f����{)쌳�bS�^4�R��ER�;Q�m�3N�#\���垞ܻ�7�Օ��3��D�_�����G��*��7�!�4�=���=���h}�a���Aj�o����Q<�GBeg�P$��J�2��0�P�?����m��K��:C������]}�m�C����e������u�?7z��h����<p��ݪp��l�F�}���1�}�g]�3
�'ɞ��wh+�p�0
B�衸5���N��H������:�%9�6O6iY~늪�R�,��D7���~]\ݟ����<������@;������&��vVt�R҈����S�T�n�<^{��A����ׅK��!��?��J�%M����6f�U@���Y�^{f�4Qg��@\����}���dg��"��qI�^$p��I�F�Ȏ߸^N�����悁>%7�o�+'��h����g���W���dE�����eݷ
�R��Ō',���w�@�.��\�	12��r!2�a�f�������)�ƒ�=��d84{T"�T��([�z8��5�L����Q���ګ��I�	R$����&���gӐbYM���������#��
�U�A"�/�q��&"�ݑ�Ί�f5CK��2�\V��	�
t���
,l��W��P.��4����6�T֪�GDKB�/h�I�A��D��w���;KWk�uJ�:�t�i�Y;�� ��6�S�#�Ǩ��NiH�sz�F���N���s�Gu��i{�u�@.L����UEx���u�6|���0.3�ԫiD��E��HR��W��,�K��ZP��[��L q�Z��T�l�L��oB�z��
R�" 2�2\'O�V�.��H��L��4�M~��L8�g%ET���
c��Z#�'��� ��p�v��9�oЃ�H�������z�}YjH#z�x��`ά�Xj;j/��Ϧ�Ҽհ�YBvT$���B�5$طV�T�Nտ+aԙdL8{��� #��?-\X!A}��ٰ��r��;��$w�	�L �;ۋ<=�t_Pn��֒u^@�������	~�R5��-?�p�C���7�v,б5mJ�7�J8����8Y�+�ܐ�#6��Եn�5�?���uҼ #��Zϯi6wk?�̥�� �3������֔N�w�$�h��k�36�����հ�: ~��fO��� ,(�}�<��w�mN���ԜA��,��� �ExG1q����P�^|���zDt�ly�R����h-���p�^�*B������C�(���
�UF*��[3���(�6���* ߩ{������)K��	Rh�C����� �}o�F������@����{��2�B^��z:k��Nn�3,��_��ʴ�^�h���*��N3��яt�rY�l��Hn�G��x���V	$`Wy�<_�EzT��]��Ԧs?0 �:�QOw�4,�i���r�0qȔ=A�%�y�p�(J9�r��,���I�d�+��l,��,��B����A�T.A�A��p�֦#O0�9n����x;zZ�_޼����!a�	͵g��oi�)�����+~�r�O�����YU�k�>��浩�C���7��7��W+�ޑ�a.�HA}
���s�0�V��%[�W�|hݲޚ�߸�NfFp����F�=��	t�&q9���f���	��}�e�1|�
.~hW�I����8��x`����-R��&'A�3$���ݬ�W��/�*��%����~�p-�\`�
꒿�}w��~���(�ڞ�lԂ�!)D �9�JE�o���b�0��!�w=�$e�ܞ���aP� �;�vnߗ�����.��j��}�5ݯ�C�Sg[� ~i-!0!%�{%|�Y�q�_�z����r�wCN�3v��n'�Ɲ��G	����Q�-���'A���\NnB6;ڴ�	O� i<@fн:��sPP�t�0'<'�j8x����':]7�s���٨�rKiH%� t�i�6�׏�;�r��A���"�(s�D�B�d��2D�Ѱ2}x,fH����0'�	��>��-D�&�i��������ɐrY��ϥ�ł��e��j�(��d��e� 	oᲣ��[�dg������Bݠ������d|Q0�p��C���Gp�����Jcn��нݯ&�{���ȼ�
�*;�Z�2ip���x�p ��J�����o��ܖMJ�OjEy.L؋[�Q�tg��KE>��y���9�mT_f��V�,Xm1EG
�����䛽/@�\����s�&�2մo��h���*��fr��;�C�!�x�酌�ĖahR���M_BY�MHѝУҒ$����d�
�/���n8�&�H��H�f��wJHx#��C$��t���k�(H�6�#�z���W��3�p��%d�@M-�Wٸ�
Q��v8�1n�ژ��8��v���3Slؐ����m�gR��{�I�G�����;��@�~�<i^E(c\��BS��v�\�)�;�:b�GW����LL���s�v[u�־��U.�pB����!PO�ϖ����(`���MΆ��)���Q=������D%�a�w�j�V�J�̋�p�S6�D2�-E_���*HE��{A9�`Is�	�����~���S�S؉_�sv�� �f�顭�G!YLpQ2_ٰ�N^��Hr�n1��[8�߅t��;eǔy�xo��	��.$�i���\ae�_���֗H���$_��~;N�,K�8l��S��y������&��ؙ����ggRٶM#��CD��F멾u���C��A-��7�Z���.��04��A
��r�6��	Yd�̌q��I���S����~PY��\��uƃ�缙�����72֩G}���QƂ>t�_�/xE�e����=�ρG�/�w���;�����DIU�+�/�k֜Ï�������a�\]�i T$/�B�����wࢄ\k�:�����{�޼����V�G��W%�q�y�;A�@Ho��Y�$[V<=+�Ok6��й�w���h���Bl�d?k�,x����"X1Lq���YL�*�\�X�Dpg��/~<�����TQ�Ζ�(�碢�3Q!�Ĺ���,C�~Wo	]���&�A(�٢��A��~Z��I��%�ݪJ�	{��A[�p�y�W1|�<����ҟ2�!Ð(�S�x�.��1��1Y��(�G�iO]�&�~���妀�������˟�`��Nj=��k1x��}/���L*���d(M�Վo��4�g�k�ZL�]k�����*kA��f���Mz�E��	��0���0�H͔�Ϧ�Q���Ad�a6���p�ZH��QﭺOQ>���0��~�OG�	��Ő���*6kl�76GpN:M|���Kh���Y������F�҄���Ӊ7��[gi��A3��ϐ�F���+k��eD�C˴i%!Y��j��eT1��������c�j����L�9,����������]C�w��ƫ2wK������5,a-y����S�qs|>��������i� Vy��`�<�����p,�fD�h/�g��Ղdw������o(��{����#^�"w�'�-l��U����&�[wM��]3�~�p�����<�K��8I"���a�t$��u����	��IH*�E:��y^���9�6n?|�&O`=�(_��e�/�y��_��x��5�`���l�7UA}͊��CQp�4c������Z,���7?�<2�&2Iy9�
������n���Acc�Ew�,�}حVo^o-�\�.d���۶� 	�v�G�raXc1u���T��F���^�Ԟ~s7�=��j31��Ǯ˞��wOە	���� ��,�h�]���*�3���+#���O�[�ܵ=d&�{�KP�=$ �ʕ|��k9X��W(a&�.����?ڕ]�=TB؏��'i����Y�>��, 6&��R��{Ԓo63�i�����las6���ʭ꾌ƟZG$�a�x�W(��o�be�Q��*o<O2�a�B�T$7�7�\���k�Utz�B0��Y��WcN���Ԋ�,\���'�<û��Q�Ƌ?9f��C�����,/Oy1��KskyI	�e�_7�j��Ek��5�^6�_�v�2�)��zV+o�t�M�o��ߟ���������I/}�h��|M��I�[d�f�Ŗ��{ѓ�Ajbk�3�1��n�"˥�r��u�@^�.���R�1��`g\��L�=?c�b
c�d@y���Q�M���FI��b�\ 	���%&Š���
�c�.҇��2�����.��f;R��e�����$�*��MLM�r�koz�Bg���~)Z���Z�5q�'t��7�>�9�z�W�4�H�fc@�,�bl�	�܊���Ak�-^LGY����� Qb)bE�TP���Š�Qh���a�n����D�ނP�z�-���i��s�~�<���}�;&d��Wf5˶�
X,�\��b݆��$�㣣�#%�u�:���b�8���7�ނ���?�P^�<`��;���f�G�&`�p�(v���&��&��apU�Z�g##M��ex<���=�&���b�G0+?�4�<B�^���i��[���	�Z.�o�1J�<�x��M��q�G�c��<�HBʻ q��	�G���^J��q���l�]W�_<���RK�������%Xy�h��%�A�}ٱ��׵���?������im�vN�+s�����c�Tꌐ%��Y�ρWR[�#�>n�w�>�^ɲ4y{ŏ��O�	dH������93�g��$�j���aC˫�W���ӂ�;��K�/���݊W�G��b��lI ^�X-�mL� �p��m��ͥa�ʓ���+aYq"�&�v�����@�.&ܳ�7�^��V�bӑ)7��?&��W���u�#���ؾ!$���4��
]HuKϯ�T�ZI������Jw�4�=eip�A���ɱV�I��0�4��S1v64�S1�|R���Qa�MG�ʶ�fɠ,G�FU��\��K���Nn�7���Y��u��j�/����2<�[AB��d/8t�Ύ�e�"ܸ�p�b}����q�~R��m �.SiL�+�=e\𧔤��;O�|�g��*R�eM\�Z{�����34����Ino����H(�-^�����e��ۇ�Bc�u@����������[�pRʅZ��>�=dG^�^��T1���De�-��1�;�Y�Ծ.�f�򗏋r�`�	2��.� k�ɜ�� N�Q8ʹٲQ�ޮ��ħz:�ܶY���UD ���`��,��:��u}�hP �3��&���u4�QA�zo�^���F���5�����O����u�=bV5�*�7��x�f��8���!M�*Լ�_��Z�.�*�F9ps��q��My���%Tq��퓖j�r�"��Y�ȴ��q��A;�쁉�T��A��G��FT�薼��Mzh��i?�����c7v��EV���K��y����(��,��,���R�I#�xE�ˮs٣2���=�eg� +�5�記�7�2��e�p�A3�8
�R��T>�늕� ]lY��jƱ�ˈ^̮5A�a�_A����Ƞ�@-���J���]G�w{�[�=nLtE��L](�}��Z2"���ݲ��h,({�-V��u{Xc�u $+K���G����a.���I��z���@DO:���j�+`gC��D~R�4���R1��8�%C\0e��㣕�Pel=���ΰ��ٍҩ��Y�����f��f�OzJ��bg�O]��T���T5"#�R~�բ�:Q]������I�6mƖd��P?�����^�
'r��&V�2_�ܡ���W��I�\s>= I}*�C��;U�]��Tf�;R������cZ1A�����[4�y�kκw/<xAv��"+�w�9~������!�sw(�˷e��O�8�ؙ��s���v���VV�����`����	�x����-�����)���|�3|D�'�����@�N$���-?j@�O�LnH�(Ś60wo�*�.s�]���`����<+�:6�w�S@#X���)ͣjq]�_Ҿ����a����m�T� ��v�ʄ�t�W�͊^����ʺ�m3�����Y���Ƌ�����>�g� �j89��ڢH_��U��)9��E���.f����#/$Q����p;Q�Ûf8�rQ�3J h�Q���	���dr���q߱�;���0d��J�*����}N�V����Dk��_�7I�/��jAl�N0���F\*x�R���=n���c���e�]0y���^muɄ�u�Sp�{U�gQ�����+�=��|xj��Z#յ���M��k���:=���z�Yd_��h�C�Uw���qQIW���<Y���d�&����{0�M	)��W"8�1����r\���I��{������ dZڏ���J���U���(��]Cs�<4qF/өi(n�5;�(�;����-ߴ����XRrǌf�Wn6��gP��vطfԎA l}�M��
�D3�au�ؗ�ԋ����d��p]���+ �	��,:O�
��Ļ���B��Cf�`~E�lIS��ؠ�>��t�e�Sl}(���JF��HpPvn��M��̕����Q�J���#��I4^��\��f1=����q�2^,b�����^Ѩ��O$�۶��]/m�*]הS`�t;[�s)[��ۭ���M8�ʿ-k^k��Ę��|�Ԧ�� �Y��nn�dF
Ȣ����pG�DN�0.�������5��c@��^��B0 Xr~z�^��
j��"�#�X5Aq���:��t!�aSa��iĎ�X��]1��S�U�Q1��|�'G��+k)H.��� ��V9��V'9	@@��R]\^Jo�$����W���v�������R�����?[��/�DW-;�� ����g�/������Ї[�<2N��N��v"��_�o�yC��6�o���TH�^χ��XdM���ˠ���S"�C����b��gx;M!	��A[���X�[H���bW�!��Wq~<��۲[�Q��'����nض���y�"��# Y����h�*�2'D)��3��MsBeW�"J�f�L5���X�L�ca��|أ��1m�> ��t���-���p�3�(��C��N�ȳ���ӁF��H�X �P�[�+Nƫ�#}��
'�P0�J�� ��`o�3������Vj���r��)���0�r�Sg7��\�&���iz�X�R��a]�+PG�v���Ԛ�����X����<��Q�2���c��D�·D�u�M�Ĥ�.�E'{m׎���^�?��c�B0py�Y�k.�zR��x����rS�~�����0^�WqT���K�].���K�Ql݈��
�J��Ե�-�gl92v��ܶ�
j��������\2�RD��]��\���)�or<�Ԭ�.��`@ś����2O�PF��e���n�;����"�h|�\�o7D�f�0����+s�uf\w���]a�(tAf�2%�T�l�Y�O#�l\�}�����W���30�=�E\���m:��&��0�c�D��B�nG�t��^
��Atr�q�x�6w�|2��C2�����As���t`�� +JRVb�%�z1zt�a8��z,T)23�K}���MO�-_�!�Qb/�^�Z)R�W�矰�|����Z� "��:1�ꙛ׺�����M��Ȳ�Eיj�x�<~��};C�Ev#��� �>�BS�G�?�#,�L���U����}�-���|�����h�4��2{�u�6���������`����k�s��?��H��& [ya�8�|�c�f�l�������$��E��TF6�$����#�4��8�jw-�0*Vi�?5?�j1�e�O���*F7O�5�8��o�*�]h�h�2w���zY�_Wl�1*�sׅ;�"���a�nF��1�ݟ�z4!.b?[1�$���I�y�wjV�P�2n
Os�ȉ%|G���1X��Y��<>���y���nX�,pGъ:jme�/��`/�p�D`�������F��Ā۾xߠ�QU�����<�N�w��*`}�:\���9�`�$Y��=׀y�1:O��������|�\�OG��m.�JS��0�Ѹ�u�Y���9!+\/�uO�ܝG���,k��=$u�&�0��_¯����4�'�?<�,�@Zՙ�&�ʼEN/�\\�lxtM�E��V���+|��5BHD���$��\Ȍ����V�^��v6�E��V��N��`���uE8��C�'z'Օ�&����^�3�`�ș��4^:����΅��L���m���5��Io l�/V-(�M'�a//*�D�z�D8yTfr_;�s�����Դ\eac����*`3����H9�����V�F_{����,�PE�w�u�˞���]	���hG�R!,- M�)~(�B<Jn�kk$���]4C}��Ëj��;�Y����%��6fƟ��i5�Y�΍/X���ZDe���<A��F��m:����./
%$g���z�Ab>����%Q��q]�FH�+M�f�$|� 0��,��	��\K�?���Lf���u=,:g۪�q�\�?���^�۷_��K=Q�{qW���2OF��&��4�_Py�Ŵu\S�>X�A*:���Wke�0PNޭ׶6Kv��t�(kj$�b�(w��ٯ�{�_/V6��I��ڙ��ȧqѩ�9^Z��Ti-.9��lH�?2�_Z�񐁩?�����bT<́i{��G�Į7qA�A�WR�M�}��L�S�y���Q���	�l�>��D\���# ���HK�i<^���P�
�4������ݘC�a~��.ƒ�p�w>G3D�ik���	��:�#p@8��	u���b{��w��E�e�
sI�7���O%E���"�9���Xm2}��X�ށ�bo�N��6�E�O�����;��aƮ8h�!�(켧l�9SJF����8�I⹑�+4w��jd��`x&�����Щĥry���&w���� ��"Kk=���hfQ�L���03 !�u��H�oϓ�}pj�4���M��	�������o�[jC�2$��4�w�CZ�t2�,���9~R]��Э�|!]�T�f�1=��&�e�Asw�jQ�.C�콷n�Ym[�K4��>���9 ꃅ�:��ck�)0�˳�?����/�1��ߋ�)�Ч�ǭ�����茎������q�>����KJ{1S뮤�K��j�����ji�-�1x����D���1��f�D�{�lQ��� WD�f�zS[��y�^��w�����p��F�|�^�]��Ph*�^�bs:���A�OZq��?��L|�ѥ� ]AQg�1Q$�c�#��=}�Ӈʋّ��J��@K��s�|��f�F�R;=}�:;s�Ͱ��i��$��+�r]1�~��"3,�L1�ZAe�ﰞ��%\Sb=�:��P�v@0��o��f�uZ/��/��TA} 
%ҶǊ�
�e��ԕK�@ >[J�RǭW�,r�5�77+�7�'���	Ϗ.��[������M �-�����gI;�Ϸ.���w���Sb!{}��b���� $�`ڵ�ڜ�6�W6рs�zh���Uun5����K�SZC���|�4ߍ����^l;��a?s$� >��z��	1N��y�ݓ�R7��F��[p�[cG���<7�Ƀ��Z�c�<���5�(GRۖ���A���A�9�K�*�:岞Y=�ؼ�'̜ݧ����(��Z����K��Z�uM#rV̷�w8+KzD]��P:�n�[d����;�\g��cK�}W@��x%�6@�Y!l� ��_Ug����<5ȳ�׍C�D;�Y?�6�MS��U�_�{���� 6Q�ǲ\s�p]e�v7Q��ֵ�������~�{�t��!� ��z���B}P����z�?k[|��
�y���F�z��ŧ&�̻�ZWz��X�X���lX��%��e֫��9e���������h�����搚�ž�r7�Ý:��Pr��CM,� �yV�VPt�Ie�/��|ne�h�"�����ڮ\��4�z��OJ`I��f;f�Y���,��_Jؾr@�`ꃟ�-���4
�D e+=�_�{������)Ո;"�d���ҥ{���qі��3���2Z;/[+�+ӑR�i�42\�x�����'wo�'��"˕��Isb�(���	�Rk�	[��r���/<������5��,�C�EN�
d���=r�22T|62I�A+F�!zه�yd�����T`|�l�75���a�w�&*�xKVׯC:7��cڄ�H�z������w���]D�!cR;R+6����)��ʌ�ɞ�O��uO�ZW������%oܹ�%�`��>�0q�o���3"c8�70�� �ij3��{�I�.�cZ���d-���}��خg<����V�x:b롖��`hD��bD՟�MzԎEp7eN`�,b�.$<nq.�v ���l���P*���5#�\4㩝Yn s@�^z��,5�nU'��8�1�Qz�,��;���A�*�x&H�TUTͶv��?�ʳv:��}Ɩm$,�P�X����6� ��XN������S�{�>Gs�kg�:]��Jw�9$�o�_C��\
\�!(8����S�� iUX324���2���~	zm�����m�d�� 
��/b�t\��OPs#q���R��r��O]A_����E6�h`ϗ��ˢ��a2D�&:�;\���� p��:���f�.����2�|c�g��y������je�Ͷ���3�D=@��ɇ�����3�e�#n���D��x�p-�
�L>kq���g��-n��
n��"�:ԛ7(c�c)�̋ƙ o`����lr͆�m3�b@����D�^hL���y�-j|kzA��UN�E���/Ǉ�5�_T��<��ܟ�4����sV�R�/��zB}4��:m_M��T�O����\�J`M���wg�u5�~A��U�0����s���?�R]s�d����{��p!�/�$E_�c���{�E��C-d�����N�e�$ap	�5T��Q�r��P"g�ZA�4ç�0�Qڛ<��z�臐��)��k���]�����f���T�z�92�p��ub����
�/�+��G���׹�b.~������o閅!���<kN�>0]�sKU:u&_���sF��|)��T��L�sV�Kj@�J�_`!��Σ�����G�,�>F�
.�~I��|v�â~���O�ʜ�?������1��7�TV�*+�� �)hj��Y����?�>)a�E: ��ܛ�'�h~u��ˀ�)�o��T���AՇ�/�5{��p3� u���L)'�z��$�4�4���R]���Hۆ�X>})F�R��]oR��/�d��T�׏�zs��k~�'����L}]��Jq,�3�N$d|�л��a�������@�8p��
�������j�P����Y/Ә��9��V��EP�����r� �R��R�@��[CTD��N^E.��!���㕡�����pJ;��;[:ў~i;S
%���/i�4���t���(�yI�/b��r����E@�,�CbTK�IT{��Ɔ�'{pz��:���p���g�h�^�٩�y�*�������!���X�K�Wؐ�^W����K��!�����:ӟb�&�$����� ���a�⻌(�n���{F�s+�elW2��]��4��u�����Ұ��<�P�����  �Z٣Hs-������A���]�x�����J�Y���n��`���iQ[}�]*��z�7��2�Qp�ķ��=�q�t�Ht��9�/��v������(e�X
JA��P��fj�u�\j��/���g���H+AuT3dk/�L�t�4'u���������"��л��'g_}����M8)�pe�F5�����#ֱ:V;3�KGK?ٶO�g���9cs9���	�膎�3\ՕȮn�Թٍ��˶?�ȴ��g̲$�SA����-^`���j��U���@�����KԢ�g�p�q�w��h��ɿJx�_ہ�to�j�%�!H֐5���E����{�.�٥�f��^��T|� (�)��U����"FA�8i$��:�d�{%���f�P�("��2/����$����p�8�^��4m�v9R���檪��j�[_�~��Г�~ؾl�'�Z>f.463GӁy1)��o���p�ch�����?#�ō�#?G�w�=B�h��~S�UH.µ�T�Nj���u��^J*{crN��
#���=��&j�����	�T-��^	�~"S.|��?�S"�5)l5hsȻ��n�LV�"B�9�^���w��0�p@X�L����L�������S�x��w�ºY2v�<G��i�^ñ�H��(K��~G�d���a��W򽲺���Xֲ�ؤ�.P1տ'���Vuf�y�+��s>y(}ơɀ�I/O���e������承��Ѕz�}�U�`ܹ��{�����/�|ַ'�j�"���K�� �BI��
C�j�*>pf�P�9d����@�oOR��=��v%�s";@ٔua�4�_T�G�%d����iٳ��;;�$SK�2kwi���o6���^��s���_PT)��la��Dȥsd����}R�-++%�+ޘK�7�I�VnQϞ���>bP}&�5;�	9v�h�wO�d�$~��xg$� ��������I��*^=�Mw�v�T�ex�?�d�4rL�iǂ��I��?
�2G��#|�d���S$�ki�r�!�Bs��2�1J[#�O�/�'8hbx�|K%O�23K�����_U������(+^����Z�U��S�Hn�-Gl6�^<>�1��W5�}p�ރ��K������"�WhA������9C���0��/v�h��X
po�U�p-��j7a6��z�=����?!Xy��ivyV3c��P����H�L��.�)���[�Y������L�W:���h1��-t�e���O؏9k��lp�6I�g[�_R\�G5�ն&����Ż�9�Ӆ����t�ٶ� �V������7>b��%=Dܑ)g���븬�iޢqʓ��kӜ}��J�r��H��$���[��-+Ks�ތV#�o�����|#]���?q{��������E�r�,-�M�vv� r`_2���ƩQ+I$n\����4��{1=K�Ԃ���D��\�7�����(m��ܝ>X�7u�����^��.|�,���#x�v-�)���&x���8;�t�B�ɮ?�=s���:�`�qV����T�\}���V����VvG��BMO����}h�R'�-+}9n@�R�lY8��]	Vh�3#f�0����aż���vY�JJ@�C�
u�Q�p����֭��
��wS�[1�������b ޢđQ&ë��v͒zhjH�N�t^ִ�Қ�x�;"2�E�jP+Dg�4"lܪ�';pZԉ9/פ4���;�HE/� "8�oݭjf��1�cP0�l����-�3|5Wit��Aܟ1��\���y���P�Ѕ2����1�r{"X��Ľ��D�=ZҶ����&UD�nQ���;C�6"V��UY��ۓ�L���4y���_<����~�H��U��;s��6�@�*s[����l�����"�? ��rO]x�	�{�����.�s�E|�,x�f�M�K��Hzӹ�w��7����V�x@ic�f���$�4�2��-�=ۭp�6���@׹��V�g��?�-p?����q��ƚXMkrE��_kC����p␫�4:�˛W�P�݇�8��0(�w�P �����=���-rd�����=.����dpfr���toř@҅�(�l�~���-�X`��9�ࣾ�Q���G��3�}��-�S��W��EHu��u< ��6�-���m�Q��}��z�4p9XyP`�&S�w�b�2�e��^YQ��T5�����Ҿ�C�X(4D;�o���/��Wq{������:�x�?��d���t�ے+�L�9���=P��*�X�hmH�Zq��M���{�A��e�א�����\���R�p�<�48�M%O�aN��ļ$H\��&��ɟ�L��h�F:,F�a44��?Q�Wb�}/8��+�P�G_B���e�F������L�N�	����fc���������ל
N�g�/<�t����:he����Kǹh������bf�Y80�4��<Yu,.zJ�qy�q��H��~f���8v�ѓ~|I��#�6������<��+u�/�����)�=[G���,`0]�Є�U��XنS� U��3`�v6X��]��?�fk���L
<��z��t��E-+�7^��~�i�r�~��W~�3^U;Y�;��[0�s��8"�3c��Y��8�|T7����X.�E+4O����r���SK��Y�����_�й,=h��@�Ы�9�n�uP�21>�*�65+�6ׄW��e��K��Vx����� �W�+�m:�����[,c�g%4q{�l:�P��
ټ1�<����2�R��璫N|o"j�/H�7��x1�U��$ȉ4` �B�;^9uo�@6@�����__Q�m��"ʬh_�7��|	c-L��l���v}�*����i��j��^�0G~�\Dkm�O�\_m�q����jjR5�L!��5(C�{�Af�~��}FGerҒ�+�)t^�\�`E�XCһ Q����y�,ԣ/v����h�yǴ�Z�׹;�p���2�sv�^�������trԠ-�����<;��|�-�S�3g�#�E���y[İYć���۽_��r�9TSo��O�ׂ&zQZ��"�"ժ4�6�	�;�ރ�f!ìe+'�/��Y�#�[3�w��������qG��Lu�5�4$�!���,��~4��{�L�Ҋ�`
� kO5������aE 7���w��G���م�}]J�?k�Aƥ��\ԬN��3��!��JB�6�I��,a��!rDݍ
������Vm��(I*Ì�c����j�V�η��%�ΣC�0B��������o��.�n�*c�F����g2>MU��1��9z)�ڷ^��yT���"�vG]tS�Խ�|�#��'��{�"�~{K�S���l�����J�� L1ш
�T%���W�j��9�#��������%&��)(�f���{��ƅ��(
b~�@3�f�)d4����Tl�w9X�ຏb��H����ԓi|r�UgtGq�҂�ow�)���+�2i��[�����AMbʐ#�8V@��Aq�36��}H����Gx�,m¶jא�2����A�]���uv�0�Ո%����:5�F9�oų�����9�JG�R�+ۙr��/��e�� Xp���\��J���k��	��Q�a`<��䢹*�a���mM y܀���jGC���}�X� i�
��E��? b,V6��Tc`�X#:���O;��_�c��j�e����:!IuK�c�'�M,��\��,,0qǺ?� e$_��Tt¢�{;*����LG��~w�&�!oR��z�W�*r�+Tk���]�s.���OJ���!�_�΍TX�E
������j����+?���Q���P����/3-3mhY#�*�Pb�ڪGy)�����`|��y�\|3��V��Ɋ�ߨm��x�sz�P)���I/���<�3�W؟;RZ3Kz�}��J�@�`�R��_��V�I��P]6���a.4y?�� �G괍�;9xu/��g?M�����k�XWB���}�Mh��c���[a�ͥK��n�˗ҫU�����6���O~���{�,E�tٺ��z���V��M��I�P[�ֽ��1]������i��y-�p>���qYp���o+9ڻ]*i�oe�M<�����������Z%�Ə�R%[;Y��d~(S�ʊ��L$86�cߊ�	]�D�D�����r��/�u~q KE����!#��6p�u��C�xM,����X��~ְ�T����e9�3>-��Yi��ȷ}�1�m�f�pNu^�ߌ��6@��c��E�>��?D �ͳ~�a�Ѭ{��qN�ښ��yЍ�8��^=ew��m�����r}�^8�~��ʷ���g���U�vyl���z�×+,1ձ4.�k�y����n�4e4�hcWd|�Q]ͅ����2�S.��%�xy�rk�p!/�hk�H�ե:v���ݫ��/�����r]��yn1��ͺ;k���/A��.�n����H��>u�	����da�T�Tf.��A�D�l"7�0 nW�}w�ا"g3�W�h�5�YXC��;f@=bC��.�����%ғ#���p辨�Cgs�Jy�;ccZk>�ݹ���������0��Ϥ�� 9�r�:~=~���ș�۲�P�<�G��F.K�%l����;6*��X�n�<��ӼDq2�q�%��ma]���/N1�˸�����tFh��- 4���v	���n�h�ڡj�*@ J�iO�������y�uwFΣ�!=V�"�i����V�c�:9tT��3�fu Ze�s��o8����1rf@1����	���]�!������M2֚d�%O����ؽp%�������I���+���j>��A2~aǥ;k�d����s[]H�eB��S��2T��#��O���2��ʠ�%R���՛���06��e���ڼ	��gW�"4�A�)�L�>���GнD�_F�����m�~܄����\>ggE5R�b�g�׶|��,�Q��ó��[�6���'K2���;���dP�}���n���&�=����Ͽx*<��f�j���C���DW�kV&��&�������V#�Ŝ�Ƨ�ߓ�j�������?4�D�
%���i�:�H��ͱwI��̌��}��(��<86�qp�=��z�������yy�s����������Ih����؜�5Ts7��+�ag�5tg?�DN����z�:;��;�\��p���pg�G5NAA�[5�/c�Z�_10<�u������Y��7O�~�d�����1��e���A���kK�[�]�c����g.���B34�xa�3��j���!2b�����t޽EG��}w�L�z�׻]�#-�r)�����.k����r�ůN,�������;���>�-I^} S��5��x��9��ڴW:@sv
Ch�w}�b�D ����x�Ǎ��a��\�n^���	�Q)\r�cx���2DAǾ^����g{Gw8*�����Wsv,'�r:[��zw�����Р����t��� a��ƞ����?�[��V�Ӹ��S.$Qs�1�벍�U�UA"G_0��8��+Y���������xB���/Ϟ��+�ˍ��:��>w������Ċ�D��ٝ����˥|����6�K5|=��v��Y&e�����?o�J��͟��s��\�q�ፗ���X�R���n0V	��srr��~����/��( ��ttha�M)s���.�ݻ�)��s&%��)!$L���|�䮴�j�Z��3"n<R����$������E��`�f��t�����o�x쎛o��Z�'��>㶱�'��C�b`�������6/d�F�1�53m&A��y�L��k>S3�\�g��յqV��I�9}`&��_]�. CDz��e%�w~r(e��L����?��� Z����s�o�Pf���)&
����.�4E��������H{��v$��I�M��;�1{}3�����De��k5��F9�\h�e�r��H$�d�\V�C��صۤ�<��|g��Ե��ū��,���
�=)�����=L"��b~`�r���Eh;=!�������8'5sʕa�0�1.�%�_����d�H_ji�~�`qRs��ʚ�8���}	q�+uU|��W�����Ş��E��e-�E1�]-���#J���R�'�6o�/�����ŝ6^��K���$�_V7��P�ѣƈ�uО3���ԑlu��I|^��N��7X[���HR��!��t�2m�^�������F~��]Ж���g��~Z�M����5�����~" 5'V/w��ݟ1��\l;	I8� Ia������a�I��k]6ET?�lm>0�ҡ[%�|Ԉ��.�q�^[N��R��F5��U����H"E��<���Փt��O�]�f0���{�%���>���/{�u�0�Kq&(HƢ`�o#�!FX�L���tV���F�Z`��H������9~�hSb9o}Tv���8DA��진����:a���>*���>�E8R�����w �5}��l�U�P;+�1d�;-�wњ<#�'�t׺;vI16��4�F�y��.`���Ţ�����Y��h�7B���7��(Q�d�u}e��e��R�1�ˑ��Sn�f^���u�~}����^���le�Ϻ+�VR����ɣ��%�s�]i)�Ӧ�J0���d���or`� ��ӌ6�#��޶�pk�����cآzx?��K����*uG�{�^0L�F5=^#~�g����%�%���RO{�=�����6�g^�z���țg:zӮ4�|�'>�\���|#�@~��G���y����z���t�� ����+��U�ʾ����,�}_^hI��fAw*���d���L����^>Y������=�J����;{BJC�S��M������Vo��ˬ�k�"�#�$?6�c߈l.%Es�ю-�	�<����3Ō�i��OX�� �b̦�k�6m��΄�+كA��������yp�/�R�Č\�.u�+�������W�ޙ��7:/��3�������J��)�/�-���PP Z'W,ǫ)6Z�?!
�y��I����7XX71���1���_�,�j�ۺf�"뷓$	��=	6�s/�ow�^��Խ{%kV�93%�#�dA�QN���$.n{$��+��Y�X�BD����bؖ?6�X{'׌ٝ�@�8���Ɏ��GU% ��r���*���2Tִ��-���5��n����=��K��dϝp��[N-�	f,�YG�d����f\GyY�|��}Z����[�	�A��E~�a��m�O}����3�*����d]՜� ��;V��nɸ�IFe��C��݂\&� @�E5�}VE6{!M�'�����/v�40ޣy��[���E+�_�~P��E����L�}��1ڲ������Zڸ}ݍ��n���3 DZ�9^ƽ=k���VK��]��J�,f1Kđ�;��;��h�&��'��q��d ����9v�%���
�pj����?4G�~��#���������K�&H9P��y�,y�*��Kd��}�U)�z��7�2k%!Df���Wc�{�Y|���ͫ��G��F�b�]�����Ri�4g��]^�I	�j@��-3J���)FΙ�Y2�E�1�K;�M����:�Y�W涘�ؑmCO\;���zeu��X��?pLs�~�H��{�-{^T �s��z����j%# �&�;�����!��l78����L\b�B��B�M�g�_��J,[~Y=���̢U�S6p)K����K��_Ӷ�eX��O�ןii���-���7������&2}��K���Y.���p�$9�/��Ϯ%��E��qfC^��K���T�@�I|������_ ��y�C�rk��`X������Zե��L�k��y��HW���Bv��������fh^�ĥ�BRg�	�#ll�F;����w��֍i�F�7����^�
���jq�[��7��륙v*Q́<��ka�/ɐ�'r��=�p�l=k����*� /r��ŶÞ�,2�� ���e���U@��^�k����)̣ ���{G�|Um��]�
��
=�m��R�i8�����H���Y~��c
�H��.e�5o�$���f���*��0l��(�Y�_IH��,�i!�A��Ė�(ՀΣ�PV{>�uGe.t�.�p�e�� ��;J���$#lY������3 l����">˂�z�ێ��曟G&x�#I�N����I���G�N����#��D}3q�B���X��{/�G��VGb���ϛ�Q�u݂���w<;Av��
 ��z�V<3�� 8&j���^xV�Sf\�ڐ�����zJ6����;��+���� ��X�!^} J�;�4xy	[��Ks)�k��<��� #-`ׯ���3`�cvD��/ܗ�]~��*��X�8ſ�*aT�=6 �
�:gn�cDc*2�T������l�]Z�"�$�e����i���e����nBTnod�߀����: @����\�s���?�4�D�Lu�*�ML���v82�?��R�C;���O����Bj���hۿ��HK['�2�σBv;�m����W�A?P⒒��r>�a�k�?��9p
�6�UK���h�t�����TzM&�{a�/\_0�����%�����H�x��P�&��OM���Yne1�X��9��Ul2vCC|I.�r�n��^�7��4N6�Q
�Xo	`����m��@\Q�5�5[�U��j?�zc�"�[���V�A�Ǣ,Ⱥ^}��������L���1�.�o1[�K)~��°I���e>�9�F��Y�3���)= +u}�b�fW�cw?l�6_ ����/ӿ� �
"�]�?�R�v������	^�
��	�9�^4.�B�l���X�~;��\�N���x%������B�Q�b�m	�#�9�X��[D��֞��S�C]�6�[����}F��7�
^�~o�m��6���/�`�ce�%�oȳ*։����~�����Qp?JL�Ϗ�V�x'-r �W�xU�?^�~��D8Qp&`)'O��1}��ȷ6*r�J�����yB�P���ݎ��g*�d�4��\�����Ù���B���]F_}P��N�/.����6��
��K�f��j�
ܵ$��tzͲ����@J�fvX��Y��hYT�t_��Qu�� k�L���ӣ��	g<�JIBա���O�II�{tb�؞̜��[���4�Bo¿Z�'{*2&�A�ǐB5��P�z��ͭV�H^RakN*�I�F�<Z�CY�M��t��W�~�Onk~�|�~.���|n��Ni�6��5d�cu��v��|���VL;1	Q{��fz"H����\F�Q�P6�����Q��/��������u�?�9�L$\{�Aʢ�<$�\�=M��tk�Spd�0G���	�.����[�LՒ��8������Q˙;��?y�0�m�|��4��B�3��qgG���'����Ŷ�,�$Z̽)FYVf�/��dg�D�q8@�kn���KRB�T=�Ӟ�}���Qn|N���~��2F1b�)@�o���+��{2o�H��4Oka�)��ҷ�:!��ڄկL�b�@�8%�� ��}��+>��m�$Һ��S�H��p�Xw#�
h� ���o<���u,�`7�Ze�m���q�{��;]m>H���A4���~�0����BMy1���U95��knU�R�]L�O��������V�)��)����������̠b�"�_���-�_
U��I��P��EP��ʹ�er 	1��C��sv�����-Uk��Mk���d��ۙW�oק�[祀��Qd=���GbR@8�uZ�P�4���+�qV��Vv���lP�A&O���9}F�%j����'A|Q+�.�	�;Z�rDBc���F��SI[��I�r�^mL��^8���sw4��7�����(a���"יF��\��b�+W;�w�"���e-wF��3��0D��f�g9W�a]�y����9\uv�O����Z�Ք ����{�t+�A>�T ��J�46'��.X�[���12���g��DW�,q�Y�OI�qVh���:�������㎔ ����d_�;�'�v7�m�4����y�����M>�x|����~��������
��F`cr'M(�*+��ŷQ��!�K n���N�D�Ԣ.�'��������JA��T�G�$Aܞj(�� "�*����n�>�����l��-r`�����HGl���OƯw�6��{yG���ҋ����^B�����g����ۡ�3��h�7�R$8y�K�*K�il�����A�д�,����`�jM)@�|�K��z
��В���B�Q�������sk����n޽�k�3�
��Dep����cb��}]o��^����Y�x~5�a�ViIH�Z�\��^2��3{�t�>�fU[��^˱�b����{��a_��U�b����ʘ-�)�84��a4�����Sde��Lqw��S{=d?s=�ͳ���U��S��P]��k%�Au­�:\�ˬ;6R�l���I����.P�ة�L������cI����FF��'Ԗ������*�vܢ;P��3j�M��B��F ��I�mOq?���0�A߹WП3j�#QF�n���(ն�l�q�E���s]��!��<��6�I��$eU�l����D	�'�{win6�ao�H]o�X��]H���"#uN3���X`?6��
��9:�ڹ����1��(B��~��M�d�^�R��������%��B�d��2����3��@��Ȃ>�V݃JJ��v���8fV~���Gv"��'��O<�_8�P�ҫ9��;�u^H>�N��I+��ꂎ滬��3˱���V~	��p�h:%�|�����N?�2�5����鍊Ur.�]	͐>�I��3��j�y��s���{�3�/�V�����z���Em��m��H��o��B�)��s���KY��d>��"�d��u�����cS�(�0K�*|k�\����t*]�Kg�x�����7����7�4�v1�4Q	B�����H��|>x؂�)~���	.7�?��,�{��e��ކ7��]�u�PF�b����G۪uK9�S����)Q���ن\]g��O�2�;h ����ǘ���7�����v� ދ�])ǋ%v�
�]"Z�ΰx��f� ��� �g�Պ:-��rYa�E�,��>������'���j�I�~��Em�w��)��Ÿk
EC^���������F /Ȁ:&���h�r�CinŐ?� �����)��j
����SO�+�-�����'	=�� s����q����r�U�)�n	;��ƠH�
�a|2 Pa����-���AϬZ�N&܈[[��?�bTb�i*x�~\ga� T��Y/|�zc$��C��g����������������2tK�3l�W� W0�]pS�K(��T�!I�)�������Qs�l��<G����5b�d�`��yB;)�NM: �7}������^�6Syq.FGJB魌�%�?,����F�vT�F��0���=�a3���<Xqb��DR�� ����pl�q�ٱR�~�m�T[2-�l�)��D7[6���B�Op��v�"Vs.�6��ڽ�N<������^��K2�⋢�GJ{��e���@�pZג�
�-ʗ#�8����d��r���@q�]�}BgOq���!�r -�pu<��< ��z���#�N�.�ur�p���Z[�~a3�;3r�X��L��:W�U#��I[��ל�uW��7����{��;'���zN�闕�6s3~��WG��v���p��Wb��`�V籾ѣ�p�L��xx��` 6��A`L�/r��X�*���RJ�b��������)?=p�6�������gM�G�\MσS3����#l|[k�~���.z8 �?��-Q�'m��_	4>�/�s�Z� � ��u6n~ݱ�z����i�iq�0��{�t�lb(�ނ�E�&��;��Z�XkɌxuEV�h	e&<M,�CMm9[F	8�r�Ri��H�Vk�Xa� �YPj-(!+M_��S7�u%�@5�`��Yz�̕��=3�si26������g����d����u�b	��Reyu��7�+ZXV�Tu�фs�m!�f��0O]��7�L���������Cq��_��>���4�8*�3v�-ɮFE1+�/R���[ꐆ2�i�m�m(�
��ߑÞa���yc��&��o�K&C��-*:&1%��@�,���ʥCsݻ��q=
x:�نo��/�\�!�?�ĭ��H+N�KӃ�Rz� ����E�!��l����s�v�q��Z5�.ٴ�?s����F$��N�7�-�HM�p�T�*�^�����xp���.�/O9G[ڴ�XP���IIT��s���X����䱒u�f\	��o��أ�W'�2�S��H��v��f]�t�,7R��	x���E0�9��_��[������PK��;Q[F����n�<-g`���!,����U�w�����E���E3D�NmS�{S��[�P;%u$:::3Љ@��VV��J5���+=�]v���։�J~	��a���{�ݳ��g�d�b��P��dO�X�~�p�SP���#�&��LF�_���=ܣʑ?�Ԕ|�[�'�})%�_�V�KY����D�����{C5nm�+��X���	R��@���ݮ	~d�U^�s�?�>{K�v!��0����%����	��k�mlŤ������n{�g9?�$||��r�����/A��(�s\!��K����#c�v�P��Z��(o-{��V�5��*1�������!o�(�I�T������W�8�&=_c&P��)<u�J�ݍ����� �05	������$a��Uq��� y�Ι�c�g�M�
:=7;��6CgJ	�C ��U{�U����%]��W�D)`��>�|^�F��(�k� |m�(����:�<5mpa^m��ă�1�n��ۊ�R��bS�}0'W��fZ��{������:�����O��2�	���-i���=|&RL|�����k0r'桲^���{�b����|ANe�際��|��A��<q� ��.���1
x�t�-�v}6���6wУ}���=3{���%S�ly��  |��҃U�%�bߢ��%�7'*����umlA��~t�� ��	�-�R*w��ݤ��g�}�iv��u���7ze�������y<���ڀ���֚ٲ�&�^>��I4�чN-� ޑ����YI��ұ�5�hAe���T�����P5�>�e���j���3+�>Z��4��>���oQNO�$�bG���%�/j���ÿ��	Ö�QN��X?8������*�}tj]Tv�"��;L�Uf����/?\>u����C���%-f3����^���ove��`7���o����3z����E����h���E��}�&))��m�lREm�}Է�3wx�X2�Pf��7=Ϸk?d]�H�	���;#���Sb=�ռ���?�A@��Yd��^��JM�8��Ҁ�^TD|�s����1�� ߏ���M�۝؟���K���ހ��v��}��/.���Ư썯��b�qVU�����3�T����7�h"�깂Ȓm�V���WdHZ�0��;C���u���x�%64�o�'���m��Ύ�x$Y�����q؅q }���8-�F��$6����'�<�j�l��}"OK�EM���;��ڢe�����ռJR���5��9�&q{ռ��=�E�c�!�  ���Z�ZQw���A�n�7	X@	����9PK/�;��QȻm�0��K)\3����W���A|2�	�";��p��_g�	THS����_o� ⍢k�.t�eV}M�����n��}|��^X�OM%n���KdM2c���>��t�ީT�]L�g���r��5�|��zk��D�p��<��(f�N4Qi,b'Z���J����,����(;�Mhq��ȑ�$h+�0�G�'��k���["5�l:��`{R��ۯ��X��y�7�����S�P�c�I͉��-4�b���ƹ�ȉs2"�o�څ�y����
 ��[UBM~���wO�@{)͆άG���Tx�����xN
��������_���I�C��]�
�~=d��A�[m]����]Qh�������w��,�'����t�@�t���H�j#{�ٯ�k��[�ڒ �2�h"�e�a��PG�qD�l��(�����zN)c?�:��|�T;��H3;�R,T�(g3�w[{��?^\hU��ɒ�]���ݾ��Q �z���b7��F����|5���{� l���q������~�L]��<���.	�t�/L���gj��۹�jTt6��^f��,�_�x�M�_��wXO��vx��= ����;���w��P����aP���+��:0JۑC�}t�a��h�h���Wmվ��s��{�-�{�n/����c��6Va+��E>���3$-�C��>U��p��ܠ��0#!�c��o�4iq�2MBlO#a7j��D��ɋ��!
?P���U��ޓ'JX��%��NA�B�<���#u6ǧU-mSܪu�K��ǂ|�
6�?kt�������*鬒�}W�o��uxz�����2)g�5fi�*	 ?���fK5��E��Y=��k�Tg|�*̬�</��I@!�lzch��zE�)�M�v_T�4X�
�"C�}�D6��q�dBʹ��7D�{W~	B� q���G�E~�>/ľUk��}yƊ�xBQ
B�a���n}����s����}�l\P@�䟻\q@�خ9�ފ@!=�l��=�F2����Q/2�;����p����4]}�d��To��ο��r���yɧ)��7��,w�n���?�/n �.�k0��,@��i��kkqF��t�@\.v+AE~�
�F�:R�9,��0��~"�	8{��+��!�����_$�{�`]"�#�
��Pio�]��a�+��Gߑ�󍲍�E�>>��	xjo�Z��|�@@XU�P��Iׄ,0�����߽��d,�d��Z%(I���E���$�!�� �p��@�Ŷg=����Vi���H��mv�>�N�lE���_��X��?4(�����_���$��2����S��gǽ�4�:�d�X�ъ�7B�g��r8�(�	�}�GF(�e=�F�h���_�/�s���)m��"~Sz�|�$�<�?%2@<�����e�b,=��ae:��d�q���zY<7�����=|��WK�X��{��~�jSa�L6a/����a�N�Ժi���d\��^�'�����iJ���80�����}[�H�a3p���3fȮ���8c�8�7�},���'"u��V�d9�Z�o��^^{u.��^�ӖP��Q%��������6λSR�Kr�/��E��Q|��ْ:���g_/��^����?���3�5b�K"q��$���lU�7���w	`��k�wcǤ14���]���3�+1 r�t�xQƿ�q~Z�[P���?�K�ah��6`զ-���}�O�Ό����4"��UW:�!f�Z���z�j�&�wQu�r�Q	�ƣ���&.�%��,8��Й�_�&�e�|�ִk1=lμ@�x&/�_Os������8�T�BČ:��cn�{��\d�:M�	ʕ�uj��̅ v~&_N��g�����)"��QP�x<x!k9���<Q^�w��$22B�+Yeyj�E��n�~*�D�
��S�M�1�4ҷ�I3����U��Xɾ�c-^Z����������2���8���T�V��Im\.��S�m��!��}��!yO�(v-����z|��*F����T�{W�����H�_��
7�}�Z"�v��+�ry>�H����Ǚ��/Z؜vD.Kw�~��}kP"��� ����b���t��R���0��B�$�܌X�J�&\����]Ș��@�X��z���}��:1O�$a ��Û�����7K�-��[a+������nnIj�~����N;��xȱ�~�{p?�:w�a�����5�`_	ܙ~ܱ�}�J�����ј��df�4ѹ5d�mÌ��7t�0�;�謹�%�2l�YN;��|��J��N�T�u���!������s���/��������mw���iݗ�����b�a?!x�w��p:�r^j�3ߑ�'8�1:�e@���y��������a�s�_K���*̟����x]Y�F��#}�a�݇���]��צ�Ȯ#Yڝ�m\��&r�-ܿ8�e�m	��Y*�$��Y��-W*{�d�y	��_��2`��su���>�/}F�� 6�V5 G��ݛ �8�3�Bs�#v��	j ~Z�1xC&�?�������-K����V&��+''O�!4���b⪪�R�*?5��#FFF�R'�)����]V���[��\t�
����χ�v��	RT�Aܓ��ư�H}�L�:?X@��_�_���t ܊�����~�/S8�l�Fz-�{ߞW�P��3�F�ib����p�v��Þ��6��A�WE�<Ӽ�=��C��!�ã�Ͻ���|�����|�ɜ,�{5O�%T�j��5M�z4V,$��/,�.D��3�.$G�Z,ʣ�sg���)����n��H�p�%��������hF��p_���n�Ec�R�AJ`�HF3�`�Vt_]=2x̧�+�e�U�JZ�>�o����W`<��]� ��Eʿȓ�0�QvTECu~C-Qb�DE���v�@���9�<-��2��/���Xө?PJN6S_>�F���+}����TsՂJ��]�ꖏ�Ph��CJi�����v���Wd���"+�	-�GX
���ƦyQ�v�;9�]v�	��nr���b�Ž�C����Vt��W�$�gk�UR�Ap�>�;�K�[���{?���?Ò�n+���vQ93�����:�J���s�姶Ս���4��>��'����~�jȽ�	��Ʒ�9ʚ�����F��������g8�_��~GQ%�Nm!I l	N�B�D�Y����/h|l���e����۱�X��8�`��W��8z��]��PO�xo��A^�o;F���]��8o��{�M��r" ��
�^��j(i7ij�x��.ד,����Uj(�Ĺ��������3�P�y�_CV�5=|�YqKP���+�B�4����-�J��V~�] u�ȖAd�,q�C<��#`SWBD9~�`L?8Ǫ�V��%��'=LW�|�M@�M�꾴v�M�l�͛A2���|��][����(�f
�hLЀ�5���{6"�����1��F��t#��+n
�f���̓E���{[�`0�W9�ʌ] =��4�%�<���d�L����ƃ��2�ܹ6��<� R�e��x�B��[�4�a�E����o��j����:�h��%��枤$<��)��=�=���)�~;��O5*U	r��kwP4�$?��"m�'i]��.��������B�4_�hau�Ab6�a ���3(1Ќ�X&�Z�����w;a<z����H\� �6,Sk�m��φ竷��`�Ó��#���V�*�����yt����V��e��'�0P�\	�������F��u]m*��2R��
}ΐ{�z���t��UuB�Y/���!��5I4k	����
�-�Ɩ��J���/���d�N��yA��:68l��,��ǋvWԝ�a�-��K����������|�j�}��<X��R�H3���O?��-̲���Jޣ��xW��v�hy�k�K�o=�Շ9�}����)�*�1�&l�Ÿ�����"�a�|�X<&��%�G9���s�+ 6�-�E@��gaoZ��j0��/�����5��E�����)9�Hɖ�e��\j��V�9�� E���ۑ�ܽ�6n<�ê߂�70�V��ȶ�A�Wr�V.���%f����]�U��tV���/{�+�Sa\�7�VE����� �$��y��c����A�xL�v��q�yD��J�h@Ր�&]A�`�HeR�(��#��<��R��Yϗ��>����"H�Yֺ�/`�0/�QZ!!5-����jBO>��%w�ZD��K�(��r��dJ�}d'ڣ�f�pg�~E�o�o	H-�|ض�����=S�̦��B[,���u����k��g�>�G8��.t@�l���� �C|��i.=&�����������IW*����!O�U.���E^�)�G��2��߷2RcITy��f�`��)tΫ:�W0+[���zxV��)����廊=H�U�C.3J
��i����)m(�04����g { rY͉���ڂ�u'@v��)��ğ¿�I>>x�k��ڮ�N/*�k�+���n�YQ���i��� ���#h`�Ek����>���N�r�J��F��������b0�<y[��
H|���(ַ�D��
Uݗt�G]� �厪�7OBઞ��,��	��z
�K.�\B8��
��b^��|M�Hj=n���>FC��l�!D�!��#��0"��?��O1Qa^����|V솫����#�ă]��>�������J�"'�e�{` �#̇���"�S83S|�d7%�����kwP�L�1�Uyd姖�/�9���\�1�<;�H�ϋ2z�]��gx(=����Ί>A��!�9-.9�>�$khht�"�vd�-�W9�W�E�</�g���m5�w��c���SS(=�agof0�=�|��G�4l��z>��%: {�1ꖝe�G��T�P|��	~�/��
հ'F�h耈v� ����k���4��W[c�g�(eΎ��o��On>T�8�"�W��k6���V�/50-':�t��U��>�O�����M�y���?̟+�l��oO7�J��0�2:����SN_e����fx��	�kN�P K�w�0j\�-���2�O�Y��#�X�d����}�^��ЯIC;sʶ���E������)�� Ff\O�g|���,Ԯ��f��=����zqT>��W�����-�5/�ڴ/>-��cg�%dx��4+��J��e+���[^a!��4׭�����(���s�{�����Ty䥖
ڱ�h���"����2RLm˗�4�[�~M:��;˧JZ_�`�a�H͔e�:��>��F21�[ah:U�Hj�Čn���*����ۚ7w�Ha�6�YqY6K|(��CL��r1���r�9�$�`k8����i�ûMx�<��o�@L;sl�	�T�_v������=<'4��j�)Ty�����Ɋ�-��ydg:	�^����-?:�h�z���0ju =f���jf��7v����0~��5��t��XZl��t	kQ����F���w�ʷ�9����헢���^x��s�|
v�b�O�N@�N�Z�<�������f���?H�]!���ZZA���9v�����,�Gs��ƞ+��t��Q�>|�v��}�u�y�R�PJ_'1�l9Le����BWx)Br�~-v��6���im-9,@�������Ūs�ڼr���/O��>�{�{��x[��hxL�aw���_���ƽ��, ��㕄$��L���T�3\�YO���/9��ڗc�*%���������;)ԡ�!��K���q) ��Ln$�50ā�?���u(bԋFٰ8q�r(��B�����#4�Ǝ�U��Oz!��Q��'e���慣��a�������5��.�
T?�v|�t��S+(��Ī1H��T3���s<�ۏ���|QkU� �N�a+��c�M���^0��w��n�y?���N��m},ڲ+1�/�u�@��H��
)Ap݁#ӑ��l�<��ph��U��{
����R z�x���]{�'=���&�8�X\tW�V\;�X2x1����]d�d9���I%U�9��a�[�M����[�.B��_9����h7�
�����+����J�{�A�͆q\��(��k�_�U\c�$�/0@��ͬ�c�:q����7��ܢr�����4�z�a�P���?�]�ɳ����,�3�	�|=-4���q����V�� ֭��*����7p���74by�_�+����{r�}|+�:���H�������=�aU¡�[s]������ʂ�{y?�F�B��]�w��5P3R?ɷI5O�/%���jnuV� q�u��ݝ�b�.a�M�"9��_����֧>v]�#�?�X{A�|�E�����7��RJ"E��WC�-_�*B��F��K��������N04P�	y��d����}�u�ڿ��^Um�x�U�2Z���4�}��\�t�	���JT��>O� ��ܔ(�f�y�>b�U@Im.�!�+����b�����Ч������n(}L�z��]i�D��}��A���2��5�>�PQc"���
����/Qt1���	,�t4O:�6OG6?u��噸5c�'���3=�k(�P����i�~����K�i��$�k�Q��&_H(��>�1�/����w/ m�,�$���k�Pm�|�����T�;БJ��=�G�*C7���	Z[?��|[�g2���+����3Li���P��p��_���4-��|�Wq�r�� ��G��IQ��5�^n�є��5��Sd`��)���\��h��^r�$�0���q1�z(O��L}·�$7���6�0G��r�_o��3Q�=Z�󢈎v#�"���4M��A%���z��aJ�*-�u���ˉn0Rۗ�v��#�j���_6N9V2��H�8�ܟhK�.�G��Xq���?}�K�,�h��0?���4/R��c��p6��)m󏘔ЏkM��5KD������gE�EKþ4��y��ۮ��=b:7v���2�[��'֒Z" ���c���E[G��9n�=�;�}��nb��d��]�f�A�f�f���^�O��:�~6����a����P���	D��_L��_�H<�i;(
{o�U���{�vm�4׋]�?��veg�����	kkY�GWﲖݚ!�{�n=��YO�W���Se�׳�?����A��S�#�R+E���WA���C�5)��+��q�����[��>�us����ɚ�0�K[iqZV�i�"��E_饯�V���e��-+}�N蘯���mz�Ū�ܜ�s� ������D�}S�K�?5c~Ʋ#y~�G-W�q��Hv�j�&c2j�����`2�h51��I�#��&?��;Y�yH.f[��g�8�h���1���w=��'�n��Fpz���� f��[��G{�o�����]ܫ���7�_#�n��_������m�iTӥ��6ґ��]V���%���n�#/,I�CQ���t6��XN�织�0���������q��!'i����گ��PN��R��Nv��.�\�ş�q<K7�z�ͨ�\��Al��y��<:^�6욈G|u�S�4[�i����ȗ��<�������z쉙���[K���d9���9���ْ�p�J&��
��#�]�SS����g泸���&�i��_����^lEY���g���Tz� ����Q���	���ZC������L����I��N�.�m׹��<�I����)�tT���(r��W8���c��Q��Z���A[���lDS�<�& S��M*p�9�s�[�t!�:�6���5���Z����xJj;�����>� ;�l3���,Ola��:⹘QBٓ�oU����]P�}օ�j������qI<�\S]�3*)9+�΍�S��2�[Ss���A��"�1���Ʊ.�,�ԙP1��^���b�''�HsOFѬ\y ��ӵ:wZ~����.�Ӆ��Y���ad�����x��5�̟���|)�[�HaF̬d(&�'�Δ~�؝B/�C<���
��1X%&ى����s�Pjj��^�6�-������a��}���+�i����{FÜ����)gc�d�Yj�c�_驪�� b�JOI�ů�Xq�Ƽ�����~s�G�+-\��>u�>��v�(NPjO xW.5,�K�@a�5+��G�$�����>k����1�ջԚ���͋�c�{�������U�����Z�5�NꮴJ��:O�2���)�'<�iɡ���Ւ �U����a����~�.���y�`���Pg`ۯ�}�Z��v����5�B1%��Z�ym�q���s3ݓ1�I6/�����FI^��,u#�v㫋|Qn���;$�Ǣ;Tsa�e×��e��C�y����O�hL��h���Q�	�V�U��>ٛ:�9sug*;� ��T�bD�O	��e�-}���
ȅk�����Sj+���5�D~0�?UIU�����mo�y(�s��*	�94@�X�e������	�=$ �u�?���0Zf���6�>�YH	S�(�NJ�W���n��� ^���"8e$�`�p�j�|�n�d���+�_�v�f٣�G���A�C�ȗ>�s����:'*��1���t��T�ߟT>��T��WȼVY!TY��5��+Y!$d\{˾���Y�ko�����|���T��=��9�y���:��MK�����5�ڹ,�rGj�[VS�+ђCX`t��i�V�JZi��d�
�G��g��B<�{d�G�
R��UmU�D�v�]���??ml�5�X8�9�J���KU�No�=���1��K�ڴ���l�W�d
ͬ��Qe�P0��4��\h��h���B6�Y"��'�8�����r�V	�uG�������E��8>�p�a��l�����΋�����=83R/��4�c��Kg�~Ԟ
?���ct(w�:�+����x�Y*�����"���	�T_ث���Gk.���;S��RS�j��ͷ��ɴyB��_[����#�{��e�!��k��1f�9o��N2:��Ǝ���V���=�36�`WO���5�ӣLw^�A���0#�w_�䋦c������[7�����f-3�}&;z��� 漹���V_ ��%��}T�5��^�ug�	2��|�I�/(�| ��k�)4��П�ÿ�(Q���f)Z�40��v��]���i(�)�Ùd�q�ɻ�Q������E�+Ɉ|���x!�yR�w�5_���j��b��</r8"~	���2��Ɋ&|�O�9aُ~9oۓHN��F>�Qh+"���h�ph��_H����=��(�qs�G�Z�i<����t��$����䊝I������2�y8YeY7-�~����B����ڋ{N��?=�}dk���mu^�y
����ф��e,y�=Q0�y���*!��USF�����T1���A��I������i�j������Mb|x�RMH���l5x���*[�n<�&7�a�ug%��R��Si�'��������z�ŝ�F������`.RǼ��{-6��;W�Ō���F#�0ES���u���b��ퟣ�*�.�3\�\Ħ�=�PB���s�z"f�蝕�[���O�I�O��~=W֦Y��?W5O<��ru	8�H�#�P��?��8������(V�mv�c��׹0���\�{I=��� ���/ ���"�r�4͠�2�����;OD����0@(?��J���9��S�3l�G�Ms��%[ܟ�������g�5�~hp*ƺBU}Dɧl�0�4����tK��EY�z<��y�q�d�N��L+_�Se��fs��[=Ȕ���_03����R�'�eS�g't&!�t�al��H�ji�h�a�$oq����=�md��e<#c���D��B�I��ħ���P�}�h�1�"ן�]"?w�8���e������������9)E��K`z"�����#(:�J|�}#�Oׅ�Al��G�����I�K$�<t���j�I��7�Y:\��E��h�"%39�]#V������- �P��_�e%K���=�5e���2���P�Hi>�/���"=bi�*od�!��?��6'1o��kl�M�A�"��Z�LpB>om(���,�),��wN�.:�"�fa�]��w�`���nQH���m��$g�NӮuҢ�+_[=B�8�6�'<S5p]�KE%]��.U�LaH�ϤQRČ�'T8�W>چ~a�Җ�1Nǥ�"�֛����vt�8\qy++
2^"�]:N@��O[�pVz�<W�^w]�=�&�E̼;jzm��׻i
�����ؠ�񰠒��ɽ��n������b�X].M۵�^��>�+�N��:b��U�.![�8�:��|g��w)!�y�jr��H�a����|-5y��*O~�ݯ��[����n�K�(�����x�a��bP��dN�ɐ/�"mt�V�ޖ��
K����`��*S�������fk�#��1�{<H�'dT0�	d1o;��R�S~.�P.a	�D$Q�N�v����AT{t��~�vt0K������9y���gʼ�n͗�ev�w�8�uQ,�U����Le��I�bP���>e�����>�O�3�S[8��_�*r�ļ<�p����+��H�1j��t�jη�=���p��x���TjAQn���}���.7�����p�E�v��c���^�kI��t�Xu]nr�m�&�2tY
��SB	���<�qɾOr�w��?�c�J�2{��x���Fϥ��x�u�$�jv�-ŧ%��L %�t�N�r{4�1�L�t*���KX>����g ��ǲ�}��j;�K�CK�Ī���N���g �oYB���jZ-7)�2unF��1�zV��ݼ�Ƹ�N�ju"9��W�@^ᔶS��q�8��B�ȼ�5!�cJ�.߹�x�(Br(��ϋ�MI�b�hr���7@�E%����I�G@HK_�E�9���?s��X����-�7�4�0�d'Fh��k�(�j�����<���W ;�X��S�V� ��)�*tV#��dz2cɧkJ��4=��m��\PK��t$>��]{&�/|�C��dMA�d��V�x�>���ny��� ��i[����<"o_�G���w�0�cCNMTOK������oӷ�Z�O�S�׼$��v��$���S7U����ti�QKO(�� 5��]`P{,�
4���}{-�:�R��z��Cs�w�����ӣ����9=pK�Z�i���Ku[��;!�9h�-q��U��W[�r�ѽNSŎ�iP ��/�̸C��X�뾷���S�1�����,;��3ױ�Զ�s�FޝɍU�yt���Q�z����Z@J�&�ɬ祋Ǐa��x~�(j�~,����~�c�'���w;�"zޏž��juL��m���f������:yp��^�����Q���"��ږ��:��sJ�������	p��bp����@��>��V��Z+WS
�E�>�]����ϯp�$�m:�տ��U�Y.I��
H�89w��b��q���S�t�����"�qb�po{s�->��{i�8�+i������Ё̈�0��7�����L�-���i5��Ҫb܏���_2�ū��*2�ThѝJD�N.�N�>hJ낲Ҽ! "G���CGR�ZǤ��䢦LB@����!1�� �z2�ӭ��^@���;���X�����S:m櫶;p�b�Փ�{}y�I���P��F�p�����c������IWg��v3�e�F��? �y��&�޸OU~�y�=Җ��S�"�o��a�m����i&|�m��˝�J�_��]<����N)su��zc4����8�}�W�C���
�F�-ݽ�NG�7�m��j��K��A� �|��`Ϡʛ�3Iq��,�x<�0�1&V_�q�ܻ���=mc{X;�x���Y��φEY#8�w�sT�v�F���Si�0VS��t�M姼������	�����f� L8Ċߑ��|��Y�bb���2$W��/=�����2_v���`��$F�j]�s�N�p��ým��������P���H]�~ƽ�(�(���х���j��1I��>�J.�FIÆ`��8�����e
\��Ď��T͑<�htb�D��o���	i�JA�al�b/����&2��r�-!�����E�"�M�X��D�7�oW�ߡ��H#�-[�NN����1�n%ĉd�
�L`�X��8l�ȹ�>k{�����@-�:=�����I�5j��<��R�d��u"�]k>����#�w�f�ũ��v�υa�_�pl��G�u|���lcP�{� �-�2E"'���,����� ��U���=�6K�I��5�&$�GFR��DG����O$Y�꫖��~��WMv�?]�p�>h.8�E�l��%]	#�F�kg]�e^�E����q'i�y���p��j��:��U�t�(��c-�M�"��Z^4�0)�E-Y:�X��)o�I k�M����wj^>��'Ax��M	ʷݧ�S¿�k!4M+�����o٣�F|dc!�M�s��!�_L^f��k[���-���G�g{6:����&Ri��n����ΰ)`E���OCY�69����4z�P0ݳ�]�N]�h��҅8pI�J�iH�l۽]�Η�����\�ú7��T�v�Ƶl��#:��e��M������牯ٸG.m��{v.����zћ�!�1���
��a�y=#z���y��Q����],���ۼ:�:	�rK	�y��ڠJ�'��A�-m�;;+C�VF��K_r΀��`s��]�쾳oV6:t�+�1�+�E��/KΑ�->��t2.+m���v�;��:��w�)��T?0�y��W�^�Iu&�ʕP͸��s¦�?P��ꠘt��wɼ�����Č�F$�&E=4a��� J	�9��$�̭��u4R5�6�.}-����q��0Gu�9E��U�}���F��aҪ3��J�Zۛ�"���{�@�74T�0�Dl�9�qV]���/<�����Z�P�:�>��r�D'!�Q}�Z�x�Q�P�ꤠ�jf��eR[;ü�h6+3J6xj�7�}غS����A$�mT'�t�:M)|}p�N�,�G8�+A[�aL�����Fnв�+������wP2�5���1�a�x�G���r�\�Տ�vŻ�Z�ޢsj��L)���J1Q��N�B+gZK�h����B�*�%�w�\�j�4��Ntz`��t��;�։DIH���t�˗�G��.�ݿ�8Ig�h�\c���6��q[J��_�[��]�p!�?��|�T��#����Hr� .�w�#�#_xHA��7���T�p̬���5�
",�w���/��E�tV/~i_�%��C v��ne5���0�ʹ��:j`W���ޒK٩s�!�:g��dd?�`�T�5�9kQ�W�ʊ�Q-�� l%�S}��>�=��'����=�����G�(%�oex�K����!��:�U���������zH���yd_^�/\�(��{�M)^*@)��hw���?�I�sɘ(йy�kk�Q�m).eg�s^QV�l��@Ux�^��OaC~��֕�>s��o�n�T��T�%�y��qB��
��,�S���ۺ��vcN�_k����PT�	t��7���g`W���l���Dh�'��HI������_!��u�b�{0Y��}'��|_��O�J�����s%���N�eDh���ƫ�U2���Ϝ�!5+���\��3�9�է�P��e"����r�����}�$4V:�@�(k��漃�T��h�3�*;?=�_��j�G�Tpq��t�Z����2��'\��Cz�T+�4�>����!ɭ��7��Gv&,Z�2�c��[�
's_	��7���&"BK؈�J�����
~��We�މ�w~��a�L�^��G�L|����zGΏ��kx����`c��cؾ�+�i9;|���r?�`'����IF��A�k�>�fk�ʻO��Ə�G��DK4��r\��e<��(I��,���E4���,#�����p��X_ilG@V+$����� ��i���-nt��a[h��>C�Wv?����p9��0���f,u]tƆ�ә8�9뛘��ӊI�jO�a~q��e�#'��.�D��!g���!kO��n��s�0%�:9��!�r��G���wpӞ4>3nZAS�8�*�juS{!Ջ�0��f�^W�:��w���������t�9h_^\�iA�ۆ`��jSZ�7�݁ɂ���У�AB>��51,҉��sJ�����F]�<��t��q:q���W1ͨ�g��ө�
GB&`�H�!6 ��)�c�P�z[x)�ud|���!)ӗL�G���&��e���#��L��P�=i$?gnVz�k�g� �h�������@I��뿷yTr��ҍ������e�[r�N���1_B.1�-��D؜���6�鴎� ˵7��8��c�6�p{h���PdEevb)�c03�-���Ɇ�0����;��ҷ�z�{�#:�(�^�ud���7x��0����ΰ�f)	-�?b�e���2�A����lDXD��BjIǪ�=X^�e����ܩ��/^/OUC5c�ΕO:�Z}^�Antěa�a.i6(�<��ڙ|$K�}IB�(������=�/�ͯ5���U^T&��Pb�bq�'��F�$K����.�IC�9֌��#�1w'��۪�^��h�g�]���6��⛆QQ�3��9�u��4!��;�b�(}_L�dJ;��|;y8~���-�IД�XԖP�鐭���w��f�?�m+��!���7s�:�uC�m4��|��V�˯�?py@�S�q�_��?E#��W �s����M��P������O�2� �a�8u<������M �/Z~(#�9�!_OCo��������r�BSb����-��\ߡ.V�T�f��etQ>Q����J#Q����AX��%��c�!����(8�������'7:w��\��J1t��+�?L͢�z>�����	�"G��.��\w>F}��	�]l����=�S��o��~��p�e���	���/�J@x��T6��T�����7.G�G~v��j���g)�c���0P3_B������OZ�X�X�kL�bz*ͅ�����Y�:�5+JqDR�a�Ms�:�Z�(���+��.�m�|�r�e���梌~�)��u,���)=�!滅�[����P0BB�CT���0�@Iw�R�)�ٸo��z1^A�{ch!�Qy-ݚ�ɿ��t�W��	���Ȳ�k8��PM>n� ����n%��_�7'�C�yZ�v��a*��-c��GB���ES��[-5���'�5y|�n�e��C5�1*�C*e� ���	��`��PjJ�\�E������'�\��=�wԆЛ�!����C��Db������Fn�i�����ʣO�hm�K#)D�O;����cI��ME�Y�喖�����S"�u�:�ը��a��<9l	�4|���/�e�� .ް#H�X�����p��	oX�1Qg����Vz��`Qi�I��.K����L7�"��|g�Gi�g3({���p$�"�;؍��� ���x����O��;��K����:/Q��J�@����"�ϼP��Y���_�Ux��_�B�?�q��<�MB�}�o���{��Y��d�ԧ�p=�x�a�߆(��㐕���b]mW�gwAn(��Pohe羭�9EZ
��k�9���ޫ<��O�{��mE#���׼�PrH�&��g�V�K��dI�R=#��W�b?�5�&�(�GRZ��fYZ6��?��-ПWV���c�Tõ�0&�6ߏ�u�`-��A6�#%�� ʔe��i��ӻ��/�7�=���ŭ��3�G�~���Ȗu������#�w�I\��й��!������o|��;��:;���3��}��)�D�q������k��u�k^e����X�y���6����XW�뮇�>�$.@:�՘Řn�r�nR'�I�Z66���[j�'2��@�,�.���nHr�,>�|���B�$ v�	�%ï]�� b�N՘��`��T����Т�*ڢ�b�Q��y��р�xS�.���H�PB��ɓu[,�nנ���~�I��'#�="s�g�n��Ѱk� �:��Ӡ,�"���!��JJ�3Լ��,��/'�<�\�,���\�H����m��a�'�_�F�%s���
�
�A�D��n7�X��Q0��6��2J�^����|x
�ĸ�� a��y	$��ee.���RB��������4tp��گ�ash"!��}�	��$C<�g�v@��9&�:��+�9�D�o��}��/��c�$�Zw�8���?����Y�L�����L���tR�@���	pT��K�ߊו�gw6�w!X����@
�Bs
��OK��g$�r�<Ri�T.Rq :~�91��5$�U�i���QHW�m�4n��L���w�h���g �_= *���z�Jc��ԛ�N�C��=���|���< �uC0�d��`����M�F3x,��y��VѳE��ݜ� ֩8�"&��8�3���9֗�R�茅�2�3�jTS��/�N�ݯ�\��6�#�趔T�`�@p��=�$T��[��>����_:����pv����13�%:�2U�'c<'�~�ëݧ���pmB��� �=*�_�e4��L���ImP�bµ����7!�
�O ���e�3��dD�cV�yU`�������[G�<�*x�"fޱo��i���м ��U�Щ^��R���`�����l'�V��H������}�q���L��k1n�9'�>g��9�k�L[��`"B���C�e?N8�YR^H��>f�G̲�t��+��"-�s^�Es_:��1��ꎿ�{v�8�}�p¦�+`��WnX@��\�����Hi#9%8WWG���x
R��3�8�i�ug���ܜ���T�I��3�����/�Y#�����R�!�|�M���~��&�3��Kv��	��\t�t2��I�����t��d�H#L�¾��m�,== Af<!P������~���5d#ߤOF*.�Ó�5�	��wG��n73Zn��D�:���Ti8K��Lj�$-<H"!Ѧ������n�V�L/�fr��O�6�OE�!���|�M�j�B���@־yy� P7A��a4���[m?h�Jȋ�:f3�C��#,L������WP�P AR��<��s���ⅇ���/m�=O_�F���gY2�����pR01���ԯ-x�̿�s���~�-ĸ|��]Ȫڻ,D�!8���=�'�z�%j��r~�kR�[���%~�i�$���W�A�x
�w���$a�ŵbt�"�Z��N�������+�rXnV�|	�v� ���S��e����嗍K�Q=V�yr&���?��!�� y(�����J��ˋ�'�������U��<��1�
����>�R&���r�����7�O&����������(+��̈�Г�}fr����'ﶺ����g�v��<��"
~�h$F�:p��+�MԌu��R��%Ni2,_�"�_��G�#g�D?��P�����"E	��cZ�P��$�7C⼬�15���/_5���J�����B�=,�ѧ���_�؊A;��B��2[�`��;����]٥+�
�o?4��5�c����Pf2�I�_����4�b��N<����$��K\�ډ��a�5��~U�4�:0>��Y8�������kښ��)�,>6VK`���r��଼�� �e��15���(VH�s���I��TɈ�����E��ݶn�#�.�-7�c͔Y�n��� Q���?:��T!IC�z?[��a�b�\�z�/]�-V*4�؁؊��h �j�3/L������_�4L3�Si똎q�rIP�λ����Ó��\q.[�1s��l�Ӽ��Sd���ۻ4%�\�T�t�+ߍt8d�=���w'�h8�x�(���"@�O*7N����;�2L��B=gH�D�?�m�8���e��(�jtt^GC���Z��I!�v����mS46��O�
�������&��
9�j[���$�w��5��!��h5�� ��
Z^�al��.c����A� ��ˏ�u����V��r_�> �lԨ�MY��Q����*�C�}�Brz���1DG��� ��Hu�Bw��> [��=^.*��5+~�#u�&�ng�.��2P\�j_�f�t�zb�$�q�ON�����>#��c�]�Y��@��5 ��.ARtV; �s���2髋�/ۡZ߇�����Zbo��?���>ۼ���l�A��~ְv-���)��T2 z��v%XC�JpT���jE���@�$�M�x�Hէ����1����<x��P�f�zk|���`���0
@�au��e����ْ}O�hw%�Q�35�w��d/VC%��
MӶ�VpXI��T�c<O_9_�D��	�z��&�[;���a�Bxq�:}�Z+{���Y�W~���Gw�M8(�뾥�<NC�Y����<Q�)��JB�=8� �L�)���	D�	=���-ޭ�����&�V�S�P��+��q��H��A�2������?{�e$,��F��!���e�(��}�o���{���ॕ�~>��v �9�/�v��o4�kΟ�s���G4w�/Gd�s����_Lvyh	�}w���1�M1N�Uߣ��ⵛ���Dd�N����:IE��t����܃��ʵ
���~
��C�^Ay~�[�?G�����g��#Z�Ql�<s�E?d!��>�Fk�s`
"G�S����5���3�T�Z��7&y'��x� �e��{	x�Rl�[��<�h|4i����0�W��<�x��P���iiIk�S�pߜ�e�Wyb��`���L?�b���Y�a9�K�����`
$zMr�U�7X�4��0K{s�5Wl	��n��XD֡�'|��v�ߵ�۠3�
�B$��>	���.^gk"���H��b���'�<!��'lQSk�=�Ջ;��	 Z��	~Ά�x?b
��8���J���R�;�Q�0^A����[z�{��݉�g�V��QY�e*����y_�l�.G�bF�\��Si7Y�[���&	��J�����^��6Ɖ�ot|Д��V�G�;�Xjb���#�~I�}ٕR4��I��1ѩAF��N��W��B
�k_0@�T�dKQA�� ��w�~Xs�s��3�xg�I��a�*��m9U�׽�`�����V�ʝ	�*9`� ��� 2��*�0xN� �u>7��U�j91�Y>�D,��i9�����ݏBU��X�3�ʃ� ��I�-��J.��"Q�pbl��mVBn;��TlZ��2ej�Ѐ�;�/�X؅p
����͐�_ɡp���ʱ�R��Dh�� G�<�,)8�=S�����J �تZ�j����X�SԸ����z���\���|fL�����:܁�qH̑�{�[=[,��cA ��]����2.W�\�j��q�-$=����"� ���Ŭ�V�W��:��uà'�ۗy��o}�g�pȧ��}ͰZi� K|���A����;�3U�}�/'r�냁�fU��b�gT�i� �B���*@V���L�ӆ�|�/N:gy��ˇ� Y�#�$�Q���/I��+
���wz�:�sR�6�o���<���	�dt�6�}9�]#�d��	��o����-K �22}�Ӟ�e_��eLl��Né��2B `^|�ړ6�V�(�c��-�4��t6�~l�_kqP9���3� �RKy�bF�1��Ԯ����w0Q�>]J�}�HQ�����>uS{� SF�ܩ�<A+z��o?��E5����r��DX|�������9<}����F4�mh+�xyU�<��>]���L�o���|T���;\���x�>9?1�>$$Ç�{y�������_yc���`�.������x1����pH�WMZtQ@��-�Ñ��iY1-�}Ag��U�@�n$���I�K��=��(U��/�*��0����E�߻�h��ޕ�E���������+9I榨��le H[Cb�^"@�AU��v�/�8B��B��;�f�/9�CA,�z���=��"E�w�2��YҼ.:�sY&�e��13���⃱ſ���Mj�Po;�}elgrM����`h�������J��9},�n3"�����=���W����ʨ1��7�M���ѷD4�t����w�r�X���Xl���<Ts��^2�� f}􏿄��R������~ ���ԥ��2Øi?Q��U@8���l�Y�o�����¥�蓼$��%V ��z�  � ��zY~�nGU�z��W)��$3��;-`�U��Oe���w_�)��ȓ)�~Ѕӗ3'�%dg�����V���Q��z=�&�,�\�ֶ6��KӇ@��I8����Z��;Zd@b��y�4�dνl��ɴ�ه�4HCM��=��4 ظ߮�K~]q�9P]z �L�xm)��-�-$��{�=�̊W<]ꖮP��'�֤N�
 �eh���iqW6����4q`-�����H�or��@N岥��?yJ�T��HLo�Dш�,d��(�G���F �Mom{���)�~��E��oԏo{>�tɔe�)4�y<�h{�n��${�B �	P�\�Yz6&�BB�����0��	�=�i�Y�^Z�^����}c}����t������+�{_�,F��o`D�'�� �W�]U�j΂�������_�Φ�go�V)5�M�N�|�"�ad�&Q�(��'w�GwhI2A�.��8f ^�J����|,�{W��w��J�D��zq씂��n�؈?9�x��� ��w|��P@��ޘ���}�px���c"s�L���e��Vi�����o[,&�������U?��'�Ȏ�@?#�w�iQ�t��Jz�A&�8�5�՝�m�w�<o���w�f�P�����n���R�U�7�KA����;?Ȣ� ����Zн;	��}W%��������ؠ*a�ѧ+�����x�i|� ����p�j^�2��kKZ����Uc<0a�L�p��TpA��_�X��=��rи��ć	���9$$ak5M�v��GS	��k�%T˶��?Z�n�`a��[�u����Jv��� -g���%'|U��u������Y��^�ߴ]�|�2?\�7Ѓʘ�3�$�7�����9a� (��6�S�y��Py����	0)�Ou|'@h�����_��6�2�F��9>�_<��i�Z�Y�u%�?�2π
^e�J,���' �N��om�n���N�^�F<{!�"q����d=�NwߞOm]d:^1�P�ޠF{�d߂�9�aMR�?��C�#�zv����3��iO�ӥ��89ٽ8J�!Uw�,�� ��C�2uk��y��>�qC�7��G4UUbK`�Yw��$�PL�i�6[2�}:��tg��H牙jcv^���+^�ʐ��������]\�x���{�mO�^Kb�?��)~5���p���k�L%��m�[@ӴGDG�vv�t[}ʘ�����*��<\o ������wu?n���3�����|����H�3��/є"�:�ЏpJ}%B��U���gE���A�-Q%�BF2j<sX�����SIL����\�C������ꅔu���K�r(���3{S�ka��[
h�=�ۼl�;�6[S�{��w�[�0�j ����!>���|x��ǅ�,aB�f.��� q�����o�������f�3�yp"�����>� ����Z&_�<}�纳�壄�
��i<e٤��X������k�s W��3�_��-G7�aM2�t���T��/҉i3�OZk<���Ѳ���<�`3�����'n�5��
v��Z�����ۄH�_�X�? �=-8zg�v�hqo=�B[,�~�M�\},��z����s ��}��C��Lp�7N9��S�]�V hO�<V�1�!����!3?�zD�,�VR�=�wcN5�SQ�P�'���p��|�;�/��t�q���L$�_�ks�^����T��� �t���'t���..�W�G�@dܞ,��6i�J����lm���A�����q��ɀT�id�e���G"�[����8�u3Ev@��K��T��6[�)�<s�6�JT<�A�p��| lր�8��LeM��qT��#�(�$�4�E�%=�� ~	i|9���v��Cv�p�jb��tjP�&acJ��D�"�`,��b�I٫���Q!:ݢ����
���<��4 ��w:�?QR R�Γ��'b���q����Z�L�U��)�3�N�-k��̓��Z���[�
�����O����9:@��6����_0@vp��\'9�Ѡi��7�=���+^�m>�h��2qx�����W�xY�E���C,��%+1��V].3ѣtě7B�BG�&w���?E��!�v������זl��&��U�
π�5�'��~��� ��F��僘�@c/���JY>�)� ���@�uK�����<��(�)j7
끨Q7��T9��B*Ap��&�9'\�YZ���3�c<#P[�O���o!��P�m�~�>�O3�����h+f�P�CѦ<������� u!�:եj���>�M� E��n>E{��(�ОE���X�I�UYَ
R��d�Jjٮ����a��+v����<t�	��� ����]�z���zbI�F �H����ˊ�9K.���V�Ե�[t��9�({h�����(M�ō�X9���r("�mǻx����n��{���$��Sό��O �Ώ�@m���MHO��2%:��!	֗Q!&���1��7Z�F/!/d���P�kOz�SB�|͡x�I a�g�KE���I��o�셇�b�i\�Ep>]:x��V�t��ay����(�}�~s�ȱ�鏇���{h=�'�,net�'dZ�4s�"����n��T��/h�Z�j~�rD���H���a�[�)W���s�[��0:���4rb�ʳ"x��aQ���@�Ĝ�tMAf���ă�W\R�������J9��ap5i��fd$=q|G���ˡ�	�~bpr@��wm���M�K2�6۞ylI[:�vk�^(�n��z��mC���r���-�T�e~ӕF�K{�k��r�`e�=���������t](���(K��P7%������S*���No�"$e M�ˣR����u����F��f�<�\��v��8��L���>! �<ȥ�|�f~"!��a85�w�m��7x�^��囝��G'.�ȧE�<.�P�z�&����SyS���z�CX-i��Y�*�A˾'Pf�Gy@�>���wh�^�3��f,��f����V&�U�U	�u��v�b��[I���ǜ��p��p%�����7%���!`f�@�z��㐏�Q�UG忲��$�}?�݉��8�}�kb0���'��@���*��(	}�/7���U8I#LX��hC����k�~��\}��'���|�Z�6������;O��κ��MivޝS��|qq��c6�\�G"o|`-�[$?��Ju��2+,�G����[j�2�?����*Yu�)�����k��e"�OzU�#��yJ��bh��v�T���x���H��oi�fOQ��^������h����7L,����͈���[?δ#J��ֵXn<��l�0�;[$������'�)�ߟ�38R!�ۮ�^J��J��5q�d��~<�
�ʈ���� HxSLY���cl� er�3AY9yE3}��	�b�2����D/����5"�Q�7<��j:UmwM���9ڵ:&>�!>���J�ˮ��-ޘ�o9U�J}G7o�:F�B2�=�Q}z-�y^fO��Sx��ӷ�V̋����ķ;r{�����sz=�V.A$�-I99Y�A�o��d+t)�D�B���!ql&��l�2���>)�4~��e�.ߧ��<'�2�@���~@��ՋR)�J%_�m���zT�4p�{�Na
�g�mh�,o �\X6�1V�����G�,B��_U6FO|��-�8_w�9���.�5�5���u����z����v��;��������h���D��/�=�kVb)�^�ߪ�y�,���P�|��ⱱ`L����O`f���;-���53��~͙ަ�1_'��L�\z�٘r��3�?�_��m���������j�c�����h�!.S٨=1�q�H�~v��������=�46�U�V�}̽t;�qc���s�X������_��O��O��Or�o�B(I��i��sXΟ1(u��+`�;Ň1A�琶W�LVzB��t+D6r���ɇ�Ҝ��;�*�aw&����`J��NJ^�б�
�1�dG�v���13��]�ݭ;���!���e��7p�NB	x+$�F�[��˄r��M;��j7K��ϋ��@nM�S���i���JgKL��L�\�G�t4/?��I���:~٥��gN&h�ڣ�a���#�;a!n)x�I�ו[���K�<��'F8 <s�΂��G:"���jY�3Fܬ��/�J��O�*�J�!AJ��i���w��r��f�ݩ�	��[�R��>�|��qﵶ̳�&`��ZnM(��.j;%��=Ҁ�1 ?��n7g�
��˘؛ԩ�����%'D1�����}�����D���Yf����-Zn�U����v����+DQ��w�y�"�"z��<�L�oJ���qZ|�75�;r����k�+�����T����V��[�o<Z��ɫ)N�1S4��G��E�c2���������E�N��+Vh2�s�TH�\k�����5ؐyq��U�?Q�:�c!��O��~�z����Q��82��^�
�пSBW׹���n��g(Kb��:>�#�����6�Z(�O�mk���\IV�5m��KO�"p��PɌ|��>��7Ύ�ɚոHh$ҏ�I�\�4t�e�թ܋�ecIʧl3�vs䘭�-ҏ����N)S�q���C�S|�ʢ����5�l2e ��� �	���f�r�,�����YG��<5�,�:uk�R�V���*���y�0`9�ٖ|56�<F�� �A������*�&����^�]?x�͚��s�b�7��O�Q�
�E���{�������m���I�!t-@�����ˑ�E�.��n��h���%�����H����9��r��//8Zz�TYr��V~��?��_�� �*�uȬ'JI�)7b�衮 q�������e�tO܁��oA�y���_�V����[�����|�8� ��Y��#I[i�28�K��<�����#2@94ܾ�1��d�}�^*'y�Z�TH������,�1�����~7���A^^�
�E��_y�	��Gc"��;�����Su&0�Gl��I�7�=����&�Q/�����"�}��޼.*�����BIB�a��97�����r��`1/��g
_z�Qx�4@�g��搵�H�!�R�kg>�3��lOD��x ��v���WP���I(�����jya0���ฉ��B/i��.T���4�G߿VT:P�*�<�R�R,̫�|�Dsؔ�����:�aK��M������+F��`�+��Y�H����E�A�z����Y�'����f�b�Z��*Bˑaռ�ʪ�?,~W���mK��S���#��;��bbh���( ����9��l�h���/k6�}��#�'S�G6�n�֡��zA���P[�}�1���g�����Y�4>�nQq�|u���ܫ����{1|��-����:��Q�@Qw�� "(�]�J���R�%(�-"Ұtw�H,(�H�t����������>�w�u�qv���s>q��]� u؄�M��Bw�m���Y<k��W����3H^K�?���p�
��G��ꫩ�VW�%1̢$I�����mC�����~���PD#�4�Z<��l��5_M}q��5vM/?�y����Ym+���Ӻh�&C�z5�-b��V�=��L�񰅭A�* D��{�􌔌�c�y���*y:��hȅ�uaI�tX�8�1��^�|(�Dԓ
�K^D�{��J+��U?��>��-��A���o��c2�qq]^-x�o��Y@{��rR(V�>�R�0nKj~W��pu�[ma*�W���2����Ų`8�5���!��?��l���[����/��O����� x�T���A��h�ϗ��� �B<3�c�y��s����;��E��r�ҫ��3O�~T��Nj�E��hJ��L'��W�>48-�GB�y~s�����o�S ��E6]�.��nk����w�_  ��W{����I�<�g�D���bܡ�h6�*���G�>�˱~�M��ydg�iʭ;�¡Κ�g���A� ؊g1t��V����(�g����dS��4G���l@�4��/yEmd�^@��]T�* ����+�fm�i��K�u��Dfg��&v�'oE�D]FQ�l:��m�(
"X�g}��Z~k���FD�ħ��P̚�l��&���3��4���t�d�D��8����2~�y6�C6�Nfi.�7c��� i�8�СE��l�������|���/��� @��"4~V���/�_����:�:���2��$6� E���g@�lq@PA���\��j�ʮ��1��xƏB"+��[!�@�S��Tۖ傍hw�:)˗4�5!�C3��FМ�*v���_�����N�-����Oo����k�'|�
��nŐ'q�A��+����8����n(&��fϘ����e� ��ۍ,� ���ac�"�s��9
�<�{��In��>9�	"����"��Mt��D��	��r[#�����ڂ$��դ��������b�P��AK�V	��i�q��`/Ɛ�2���.z�����������Y�Z��\2;ƥv{��ܺ+4��L�Q~M7KȩK�f-�~��&�	t�o|�%����`��E'� (C�٪�LJ��gy��pq�7��O�ǿⴿF(����4��?+�Uգ=~���֣$a�� �n���@P©ϒ����O����9�e��gˉi�z
�U|�mھ�h��eй�dN�E+�������Z. ��秅�ƸČP�D�q�il=���Z��v�a��PG�!8�32ܟ��A�	'j�K�|�˭��ϳ���I����/[����8K8˳�ᘘ<)�V593N궷�a����q�}}���+�o-m����`�ot#l�b��YgP胋��p�0��]�+�$,H���J�f֤�qH ���������GL���$�:"�0�}���C���?��I����5�[��m��" ɶ�6�Z�>p�D*�aqJ?|vȒ�ߵK�pt�݆��
�E�5x�E'��R^�9<c߃B���'�.�7낔�f�% ���C����̇�����7�dr�����Znt�	�T��a�Y�F>��E�p��vǎ�_m�W	���^i����	��\��f\U���tJG&f��"������J*>�9x��\��nRQ���k��<��U�����/e�*�/����oUޤ�hŧ�E]}��FT �0=;�\jE�o��'��7�-������V�e8���X�"� H��7o�y��}'�65�hq@Ő�Į�A�|o�R��E�p3�Q����X���r} ��{��������B�Ъ`�c��{_ʖs��vf�ټ_�xV�s'�� O��?�����;������+��_�x=���-�;-�&�O�ƨ�!BD�qnYP�w��T[7U+�5��=+ؽ���n
�5vu�ۢn!z2p+���:���]�O��������(9f�4�E<�W,�.d�>ϫ�)K�5x̭�Ƴz�R��Q&�3C�%ǌxS8K��#-&��u\J&�wu����ͳM��	��*�ć��=A��bI��o˅�6�!6`�:�<�~!�/�?�nS^�q�z��8nN�TB�)G�kL��2i����"�t�Γ")l<�H��cV׽�H�L�z)g����6)������$͌O�6��z�3R#"�"��9�y��wg��lP�dpֱb�����#�8p��)�c|Z�Lփ��P����D�@�4�Y�ѸͰ��{ZW��t5��Y���i���(UȌܗL$�'%��[��Q����9�����(���1[7��mPo-�N�$,����|��)�v7*$x.�����I?��3���_��䨗 2=^<m׿+��	~ʹy��F�,� ���ӧ�x�wA��`��:
��t��"�!�����[��-@~fA�Og�9虂Sg�fN�T*�tC��;%D%P��b=vg��z`�'A�uLnaY�
W�1�#�*�~ȫ*��k�h�f���6-ȴ62Xh����5��G����	֜u?�ʽ��? �)<30sn/�b�)!j(���u�׵^�LI��5��>?�8�q�K(�a9���Pm����Vg)���c�Ą���a��&E���~;z��L��p�Υ�%f���â�6[�c���8�����h*@��+
�Wiu�P	Iɇ��ݨ�^���$�݄��z�?�,٪B��6���X_�0r�6�Gy�k	��!F���G���Y��ر���5����Y����V+/�XÙl�V).L��h�����GHL�f> 2��r����@DK��i�����&LPS9ţ�������$��8�sI\�12e��p6I�����e!'������?�]��#;�?�E�2f;?��.��}:W�������-��DS���i�/��X�ƹ�N��h1��H>;3=�,6�FCl�z&�wxa8��ӌ@ek��<>ٍP�<���ۧ�4s/!�Y��|���%�.sfd��n�{3��>�)�'n��V�Nkqt����D�@��2hk��� YG�P:0�8(OiW���t>%�{��+JcE��@}������@7��H/
ݕ��+g��/`�%��ė��ex�C�J��� \	ܱ���"�l�Uc��zk�Y�b4(�W�:�;���^j�K���G��:@�Y���4�=��wK��;;e;kS��_i���ȴ���z�Gx�����tw��G�^t����Ond{�љ�W�A���益�ln��ɛ8�h3{?��Gu��Z�7Qע^xz|`X/�ƪW��oج0�����r�	�+�@����ʦ�B �3S��M�|̻�)�@�z��V��l6���=p�
�UC�@���z6��f��s�&p{�Z0�����5t��}�o��J^���\O�s�r���&Չ`�
1��M�a��I���K8��-����,.��_�������y3�+
�o����'b�a,�����T3Gq�w]�D��b"��*`��\)����?�yy���Wd�����
^J�Ӽ��q��/���J�3��$��y�����V��Ё0���_�N������We����/E�\�v3-�*�@�p��W��	�q�*��� 
-(f���v�z���LO�� �Weuw*�4����;E�@F1�:���Ŋ��!z�F����j$��sXk�qyA»��xɘ��S�)[���t�4�fu��?ɂ�C����cv.�{�m�K�4���`�S'`��"�IłZ�_R���*����-�Q�eb��(�?Q���k����SR�Uo.�P�����h�f��Q
�R�����L/����|m�a?�P�a�o�o'�����`�t��l�s��6��0��A�nQ�ł�K�+��B�o
�R� .FT�U��_�������~p�2�^D��G�7�� nM׫��\kʙ�u�v�V��=,y�L4Q��c�P��^e>/�/Џ�1rTC��^��$.��7�B��&DzYbk�́�Ke�s���r�ϡ��1֮88�^����Z�0�/����9ب�:�f"1��C;�@Y��d�B�}�k�?�9��������;��D&�Es�#�윂��U%6���!|��W�J��Ex_�ߵV���W�JMp�U����ݡ��<�5)�]I��NB��Ꟊ&�/6�|�x�"��R(��66d	�i�ǔ�y(N�.�����mI<�� ]�l�Y��T���
�^���]&�!o�^�H�1x��;H��&3��0�D,G��:ug4�q�
�$rM����#��{�0H� ,TC��iK�;�:�p���"��� 6��<��G2�i�w3G���p�l�t�|����Nv��p�����2<��Wm�!8�iH��4rN��L����!M�Y�r��e~w��K��`-)�)�I��J��Y�TH�j�]>D3d�S@\Y���!��|	aM��t3��O.���G�QgW���1���C�Oy]Ϭ7Ͱ/T �W?W�<jhG~J�{J�ߌ�TE�E�����AŒ�^/Z�D:��
���k���d�߿�9j�� �Q%А���^ܾ�.@Iz3NY8ш�a��SW����yǯ�gq
���������.n��<Rʇ��G��� ��V�lD}8���J19h���?O|Q��:�/�!����άVKH�n����c��a�Q�>�ʬ\�X�I5)-����:����;�;q�Dz�dgd�\�Y��wۀS�g7è���uc�g�o����4�k��o�b.T��B�$���d��o7�K7��aV�%�԰f-%�=��?ح�]XE�y���(u,��2&�+����jM���Q���K�����|��[*��\���8�� .XR�~��]���b�=y��Y	���� ��=��zkZ)�h�(sq{7�����Ku���ޘ��vl�T ����z=&9���>d���lB���o8��+z���� G�
�S������D|���"�:�C�e�74�Ɯ��j���D��4N"�R4i��y��p߮���M��G�n��*��
�/���D↭ޱ�Jca��eey8r���о24m�gi��ȍ��yѝK>�sz��.�0�iWQ*n�Y�i%��D�9�Ky'4�s0�8�&��in�w̧��#?����%�9�?O��b��`����6&�hc�Ÿ���|W�;�$G�'q<�J!]�6((
�������/N�u�ng5.�҉b�b(���J;4��2?_暆�+��5w�l+��t3#��J;�$i�N.5=T|��!����1�fD��i��� GR*��j�j!�]W��1HG3# ҕl���B�l�Z�Ǹ�}�5܅x�iL74�c~����C��-u���J�~݅]��m�1<_��1�X?Vv��,j���q�� &�W����C⣶�������X�/M�󯌝�3�73�1��M��`)�3i�WɄcF��>�]=�U�#��BY�D#�]ݿ灤<�8�:��S�� ��ǋ����9�ˑ8�;�����U/���;x1�*1��u���Z�V��PN(4��l��eJ)���@X��a�!;�<"%��<��[�1UK�Θ^k� l.�q�6�l��`j�%�K?����|��#%�|�P�43����?6%��:��e;�;�q./��;(8j���I�B���H ��gOQڔ0 �}�0l���J��͉�)5�ZM(du�Oê��b3�T�8$;�����+�}Or���o�a�a���߇gi,�]��O��?r����e��q.��g������+���y}�/��L�8\<�T9���K���|���U�;�Y���w�����ĀM"	�+�-�1A�3U�j,�jу�́���KNB�Nܺ�i3�n5���<<�#FZ ���c��3��j����f!0o�$ txF�a�Qх��������j9����d�c�N�\$�x2����_���u�ڤ����3_���PG"3�Uv"���̂��-�գu��pm/��ـ�_n�����
�����>��BNu�,*+�e�t�R���6 �<=-��^<��ƌP��M4�5��3	Jt8C"ud�}wH���W�!J6�/����H:��
�v�$�7s9~O��Rb��2��W����n�#6���5�G��Ks,���|6�|�5.$|�@PS� \!��?55�{j�XѲڸ�n��GzKP�۴����5�IA}�B_�Q��&빏G�Jw3�i� �\��~��]�8c.Ҳ�M���x�#����BKԛN�@��M�s���Th�2�v-�>M�*��Q�̓.�����4�	3TV3 A%m�a�v2G���A�k�I��U�g4"�����msw%qyq3"n�n9R�	��Ѣ���t�H���Ђ��l!�2S�T���X�e�@��Ć��Kʤ�h�*�p��e&Jy�(�Z2��x��$;������o5����4���=&��H駊�O�����g��:����V��874${��c��z�� ?m%P�n�?����8�LjE�M���r偦��].�O��t�tY�Y�|,`f�<�Tˏ�RM���H��d�ݘ���=򱥹t�^�<�IBb|��	|A��%�`��pj�(3�Ѫ����慖��w�r�	�!T�'K=������nV����l�O���s�3 ���"��u�=KL���qB�f�LJ�	
��5���g�[���/��ȵQ䣍]t2�����̻�/k��@��,NW%T���q@v��#B�+�1��jE|<��ҁ����Om]|�!R?*�hRC�	�zd���x۬��L �ʽ(AM4uu���'��&��$�2��� 'r4TW}II���5� ���xB�ߩ�������yJ�rJG�ԟ\�}:�[�*.��GS�m2����O��H��?ؽ��0�~+r��GU�����"OjC�i:�$y�3�a��߱^T��2��X���u-$|fd��&�KT�1�@F�N ZYٍ��A&���9e_2�)��\�@�'P�m3�].��1Nυ�2��P3��=�$�F{W~�a��
C!yg�u~���l�FA�JE酏TK�8���!]����eXcW�xxn`u����F�5C�C��D[�Q�pda5��5��W�2�l��޷���_8)]MV1g���|ȯJ[~D���N�����.��7����@*���]]1�̔�%\��%!��������lK�{�KP�ɷ�ٺc.��7�Iv��9��IϪ�?��7V����+1��$b��HG^E�A�/`qdN&F|ϙ�Њ��1�<�*��8��&7&�` �Q���p)�J��\i�w��r�cŰ����.���<�B��7IG�h.���b,�b�a1��-.]�����7�@X&�jb������DLPf;(&�lX�%m<N�p�,��4Hx��:Q���gH�I ���(Y�ٔܚ�>�{��2S�=��\Y#ݽ��O*<̯_p�V�-��'Կ�d빃�(5�MdWV�m0Nu��RF.բ푔�� ����� $Mz�'�i�L|���R懇 _ͷnNGQB2�By���_�7^��6�B���rrX�B�r].�8�?�x����C������-�3�{��Fk,�sI�,ޝ��D��i��D�L�M<Z��yM�L|����Y�!Q������� ���L�H_����yR�%=����:��z8n.�`��s��)>�@������xV�E B �V'�ah�)�j~f�@X5�b���/�k��Xu�0?�r�����J�nM�_�H�=3�;o��ž+��?��[��0_��т�O�k�^��@�+��fՊ�
Vj\X>V:��:�����I_y�����o6��\��A���7'2//s��mA�k[�b�����9�aBX�����5�s9�!"ƂȘ�6��f��p�s�Y3Li�D%{&�����I+pAj�nݮ���C&J�p����&��>���9��G>p���;|ֹ��-r짿 ��<�y
����gCX�-���W�����Y��B�����0$��!-oT|9,��+�Wˣ����k� Vy�w�H�Aȶ��h%�j��?���{�B�5x�QJ
^I��,xވzt�����|�I�X��7���-�d̴^�%ngCu���Ě�S�����i_��s�.�i5�ЀX����ĕ�s�g/ �F��߶�U_�rƙO��������w�	�5��<�q՛����<�D8E,V��Ǧd�S��{��YXl<aRh�����5I�^���K�f�`�ֳ���3�2W��.�?���8��_+P�1������M��f1j��B�?�UH��4����� s��S�~^���K4��=��Ѯ�1c�3��L���)���K����e�Aa���g��qZ�Ti��_�����̷)���������E��<�ȭ�K�2n�)��dĴ� _tUQ�� ����r�?���xh+��A5C��N���K�.���w|�����3�IM��^t|�F�^��WSs�q�홭����6q�i� ��Ĩ����N��sH�=��P�rD�h�����A h�2 �OӭgJ�d�MH>���j��e�Z"x���hz ��;DL����֚BC7�Y�9>���g%A��ͅf���:`'��p�\��9"
�E�]ic%K���j7�$j����Y�P�!���t��؟
�
��X-rA�o"��e <U��SHu+4�¼|�m��������n�ɣ�2���N �G��wT;����d6ku��uh9ܟ�WT�nv����L��� 
�L�u�8�U�E%Iv��||�iS�* ��E"v����v�6��j������R���; U���ܶ�pb�I� F(�����d�C�,g>�5���wݞ�,�8u~�>w�#":��L�b�Y$Ԥ<d8i�q$*D_�����h���M����1౛ICx��g^U��Q�,��8 ���̀�p��mg{|s�2��Yp �J	P�:���s_�E8��N��? ���a��0����e�4H�cz���a;~\�ϻmu�A���ݒ�g�1;P�K��B]K�͇[���՗�{���M�<{Hq3Xa�ۓ$7>���aTh��	߳3߂;�1?��٘ 
n��@4�6f��  �ө�	�������i�U�d6�M{��NMK%�}5���)ݯ�.uRk|U��yj1�j���-������˾mA��G%>d��`��k\��Bo�WY��)�9�y��fi��=��!���a5ː�?6��%u��n3��|��rf�����t�@�x�FF4�69�1�x�D�?���,��6�d3_Tl�*k5�m�g+�w}�\���K����j-��[M���{B)���M�L�V�L6���;��DP1%n�W�'� ����x��" =q�q�p�p�����B�c*z��'+:��Ϝ�d��&�;�:/=�tCI�1�I[�D��رw`E�>i�:��A Agz�K&&,���1�,99��)k�k�6�ӝF�v�Q�6<6����|��P�4td޷^�i1�Z��"`��r�ןػ�2�Ñ�8Br_B�⏷�)����T�S�X�{|�y+��zgL{�KƶE�>~�' |�65�����݋�b�����D��i�45)II�����4@a4�6���1C��#�Q�ҧ}�l�G!C��!9*�*�b#��cZM�mZ7�z�[���
.�b&������ D�#��-�\ڎF1:C�|*�P��:�x>��)�9o

���ih�����^-9"O�]Y�,Ii�'@)�W�8m�8g��f.țc���\j��0�:}�6�V��Aƞ]Q��D����;�
{�6�� q6ܹ��\à�iw�!��Ѝd�Ҹ���8��4��~��4ӽ�RJO�+$X���@1�����	�G�4��C� �P��X����4�b��>x�c�̤���y^6�ǃ:df.6?��h�6�|$�O����Pܿx���1�Yǈq��Hs�&	�䨗[�1�f�&�>���(��@y�9�ѾP�R`��Ί���%g$�G��;/�i��~Q�ڮ+<���8���,x�A�官u����PO���� �E�����́��/��ߠ�W��mY�`��΋��VU
Q�	 ��J�b����`��LFFf�V@0d�� �K8��֊��}��
���w7�y	�o���.�F��yf���'d ���E�p�6KFשYD�ڤab�,��0�/M���(�k��� �����]��^��;����D��R� �5�x��&�҅ ����Ż�8��I?>����E/�4��p�Xo}En�DȱB�݈LDMk��9�|U#���1�u9�PK�^�l0�tj���n'�07���|�`w(��{>�x.�1qy��`
��8s@�nxi�<HPD�ɠh����������E��Ia�n�y���I��P�lسSR��&�b��aW:�.bw"�1���JZ�dZf>$�$Y��	`hr���y`���gZ|�����P`G+�e~�8z�mK�'�z�Iܒ-���P�>mS��h���Y]G;:-���B,�%��+�� ~ �Yҝ@��S�ہ�H=Mb�d��(�$��+O\@��d	k�{*��D��$�3U!�λP�m��u^J��6������HcIu~c�^2��tﾈ?���FR҉mh&��) L'�4({d;�"rTy
|��?�R�C������=L�n��Y��T����� �zx�ηt�C-~�����<��z�5���6��d��׎?����G���� �˞�n��N��{�����(!%�>8�<r���."y\�H�쏰Z�/RJI9��5�h�ߦ��?����zD�k��{��<]�%4Sq9���Y��;d{���p����я>�h��oQ��i�q9kC&%\5R4x�|��,�e������Kϛ�߯DV��~�7�ܧ�/�����XB� K"� �S�=�DN���8����;�)'{n5u]<��+��٣t�Ͽ3����wa�Io���Z�
�ƻ'6����v9%���
�~V������5��ҫM���5����U&�ŤM4�U۝��y�M�Uh^�t�l 򥖀���&���*�[� o��L���O���R�//$%ٗ<���O#�\~-M������Px����N���TK jK=����-�Wr�؆����ΐ��i3!�{��|7펺i���N�\i���5�}�}�*�b1*��[	�r�{CI��W�%�,%,�*Ҭ�S������B�7�H,��@\����h +�:�oRnmA�`�/&�F�Q j  �}~M��w��Q-1�l����p�W����`�^P&y���^&r����Ԓ��$���^\�
��ƾ���o�]M����O���"��e\~���Y�^�\w�$9�y�����9(����{oe���@`� %ߣ��cW&ĴAi�9m��X1io�{����lV&��<�Hh�+򈎺"Ƚk%����o�3�����p�����V7��Z?���U� �p�8֡[�2b��ͮ���X�i�Ps��k2~�a��<��N ֣�w��L�_ш�6�qp&0�{U����A���~�mE����i�#�����!�����%�I�!#kç��mt�ٰ�-��I�1�#�ZfIt �����bگ6�L����GjQh��2�j>��$]s��P�G���P�����8S
Wm/��c��������>��o�Y�}0Ww#�KF������ Ŵ��K1@�l�a��72F\�R��'LH��<g4"���e�ǋEirʄa�����Ӗ<H�K�R��J <���c%3�������;{r}�p�5A�/�R����v%р�ڽ�x!Z,Uۨ����0󮙛�S_�d&��B����B�H���D�2�I+aL �3CA��C����<[������MJ��Ɠ(� +:ۋ�R��L�mr,H���p�n� �Ky!g��UNAݪ�e���f¤�ݎ/�>�״2�sx4dq;9�`%MT@A@��*�P�kg}��k(S�ߟJ!L�%D���3� �%1������ȹ�m�3�Jһ�N��S��%,`�υ���q�_�n�[C/c�e�c�FJ?=젥"�oˬ�B%_��Hu%�O&�k�;ւ������^���-E!�q_s7��O�.㟎�'�=ǒ�����_� ����G�����כy�V�5`y��2E6� <��h��&�R�)���C8 m�R��Ke4Yᢏq���NBbsZ�ӻ{����
�;	;E8��-��E�<q?]��2��J��UA��/��*���8��,衫�o���H�G�J?�\�af���}�lY�����A[���UB���I�r:٤������`�l_�vB���p� �-����>� «2��D��%}rO�~�%����U=Am���
��7�:vz��*��ޔ���'y\��8�����$7�jŴ�k��TjAD@B��d��S��ֵ>���������$b��ߎ�W���2K Rb�e��/�8������l�d �=�.�Sl�f>2#N�@L�1,	]������~Z��O���<�6!��.��y[wU�`$�[m_��1w�h���h3���"�T��0�h;�X�.
E����dՊ�a�O�ՍyS�ԤW�_��jC�hoPa|���o���(�=�S9P���� ,C�*�k��dj��2^-�A�����۷��l�F�q!���-�y�a/�J�;�٪[��y"ST�Zuw}TB c���w��j�&1���s�HԨ�S��:�W��j�r�: 4,u|�]?��D��@b/��o;�R(��_ׯ��7|����5���������nio�i�Y1=��f[�p\-�v��au/	�0�SL��>�+�z��tq���tw�29�|�˩�c��p�'o�Q��|�"h26#��R��1�T�����o�Au=哃�ʩ{%I�׿V����7��Է�Ќ���@7��X%{��y��D\� ��y_��aW��M���}��ݛ+�GE����c7�?���������
q��vs�0�A��F$���a��3��z�	�:n8��S��[Bj����u��ί�_[��w �烘�..X�����`h�;����8hf(\VIK!P9��Vr:11Ce��ԝ!ѕ=b���Z�#��GPs�T�I
 q)Y	��<㩫���s_���qI�3�K��ͮh�\�ĵ-�2���*"�/v���#�o�E�����O�S�g:f%rn^֭=�&/�t nl�p�  ޸"KF}��i�3TR2�]��L�&p� u��"T�P%p�4�� ���V�� d�� 8f��l��L�e��c
E����2b�I�?�/���D��?i?U˃�I>/�E�k�w Yۻ�~�C����h}|�Zt��|��O�n0�$GU�;��Z���=>?}'ۆ��� ���C�I�kZ�\궸S��Y�|U�U�b<����M�#�^ oL{waչכ!&-y6L��Ndk����:�׹���8^; �)��χ�9�Hr��3��������z¤Vl����>)��7��Aq�sa�\�L�xw����*:��/P'5�|��nߧ�~fo�@��Qɹ5[n�-5�aF������_Z<���rR��K��m��g�V�ڽU "?�(�����;6�S(F��/7ٕ�4�l�0�6>�͒헛ō���h<,�!��������MOT�mr�F�yNTÙ$_;�2PI|ک�D�g�k����
Mi������/�(���I:�P��X�W�=���4V���m��Hq2?�g�\]��%��$��#9� 5���┬Lm�p��| ��AT��zg4o�o�L	<j�~]��Hx{���w�!2�1&"Ι���䴭�nb��]:b>�O^)��x3S0p���x^�N�+%	�+����s3:�#����T�����#���;{ǔ����o3e�uо���%����4��^���#����wT;����7�����l<7Fhf;[�����A��=�9�k� ί�Ԯ2yEF��q#����I�&>rt�`a��̄���l��7"&���iE�q���y/iM�[��M�B�2��y
�VW��V�2�9a}h�Vl�wB�X�JN��s����������o�������ז�)�^[��.�7������dNbp�6A1��uW)z����r*�x)�4�\Y�^I��"a�L)���<�O$_�V��[a�-���]�.���z��������Ε�w��n�6���`�m�f	�7�'�Zʙ��!���4���'�%d����F����O�E��<����O5BZ��n!*5�,��繊 p�g�@����8���G��ę���W+��41�p���z�|~��l����M� Y	������-A�`ɟ�jjEc���^lP�V�l�">� ���me�.^����!p�R� :^�M	X�ߧ���7�Ƌ؁5&�
?����>�d���L `sl�Qox6���v���~u��=�w��a��M~��N�c���9A�6폄z�ƙr�%�>u�n������V��o�B�G��7I����m�Z���v�i.b(���ُ3��6D��˞�_��@>wٌ�!����e�<MX��� ��d��!b|����ӽ������i]Tʳ�z����4�J��Ze�R��cQ�l+��¯Xp�\�a"�h2�|�(T���q�/O��{��EΓ){��v�N��3�ym�C��_S�'c�����in�q��U������?�sO��e"�N��)T�C$�'���&9�i5)�Ե������h�\�a�s`�7�nGu7gg�k��� ��M�J;�:
=�����E����-�8uOP���~���DD���tn�~�i��;�5
�ҡ<�~����/xb�Y�m��U��Q@��v-��E�]����&�U�ٱ^}����F�L��y�񜺃=� �h7�h�+t��+���q�H�݅;�ZPHU����c�������������W2z_y�:�x��7yjex�P�u�`�>~�e#j�w�t�(x�{��!_�ׅ��T����a���G�cڷiCM��ޕ�V:V�e�8�8�$B"2��%ʆ'��B3�]��
GW4<;-?l�vlUf�}�9��bh��K��5��,�E��\.
""��b�
��!n1�$T^s���\1 �)}�'���D����ۖ�w=R�����v��MN����5)��[�����#hRH�)�F��O��(��xU�^�;������PZ@�i�5�hV���&�rs��F�O�R�F����|;�H��k�8�k-wK
6�RsJ�y��d=)���N�7��%wpk�� ���4ҏ��hM��o�u�d1P�w��O���t<�۩}ޠ�w����N4;�x��W)uDQ��zLO��6��=Y^�����q��&9l��0j ��,�-3��:��ahn[�2��:��8�`C'�eY/OsÝH��lp��p�YYHH�����}]�B��sq��I��O�Sq$��iIJ�53�T�1�Q0��	i�Ҩ�o�)���\r��q���B?���1��5�0^ETw S���FEg̉~vF~�opg��"���j1�����%$n���`�,8g||w�����߲@BB�ŜEFz��U9�Hrہ��GɄ��h�v�a��޽~�1<��U�����wQ�ɐ��0l�̺2̠K.%�N�|9���掤|�4�aH�=;g�wW�s���I�ZC�Kg,�"{�o3�!{= ����p�h3�]�8i
pD7�̒G/�d�k���<��U��̋�o\���ّ�F pi��?�	��i(~�E���w�7l�T;�顫��FŒ��\��'�ƭŕu��]�����XkO�$%��/G{��>�5qo؏W��5�w1��e�(�qil�K_�[z�YPŌ-��I�����Y6�;r�(WᱜyFC����y��m:#�����iA�`�<�)x��sk��;\;�9�K"��z80�S?�V��*��`N�|q�{��Vv
�=_���	h� �Ӂ������s�J�[��+DUr�l���_�!��&�}�!J��Ea�U�]Y�ܝy�z�B��8�9I�`����y��T>�����،w����e��neֱ-p,�8�0	,L~�j��͑��	$ύ���<1��w�+��束�dN\��)�������T��(D}�Wv�G�ukBe��V���e]v��/�t�p$�3�����x T z��JI�v{�8��پa�
�����&j�)�z�����~GE�a�8�	]��r�VR�Κ�w�%sݽ��������\�oeH&�7��^���n['7���O�f�ndu�m���9Q���x��3C�E�!��$u��{[A�����9ش�.q'Q����c��^|���a��]��������iܱ{� ���H&}
 O|T�Uc��_�䡘��@����.�����[����Qmt��;T��aS\+�I��Zm�~g8{�PTLE$E@�L+�Y_�R���S5i���������uP��U,R���_�8� q��X	�?=����r���uJ�(�:�2�If��#��Q �䡻}����w��*R��=���!UYٙ��Ƞ�i:9S?D�2O�����G�7#g������W ��G��	�����1��cַwA��ǵ��Uψ<Kw���8	��ͥ��?{ƫ�߽��m�N�O�d㭘8�;��Jt��Ib��? k)��`��U"we�TN�E������u8����$�[�5V��_7UJ��g�0結"���qg�tr���b3�O㡩��h�+Ӕ�j8 ���QẏZ�f���W@E�D}/��R(a"(�"���J���(,!%,]*
J��ҹt�"- ���R²t�7�����g�g�ν��3�tS��.[�(��V�j��G~�+Xak�F�<㙪���_Wg�&t�����4��O8�`{2�i,H�\��V_^�d��O�D�5��s oH�3;����d)[ �g��FH8��+�r�q������g9�n�����sC3��0O���)3��V%�Cv�v�a��&hE�󎎇�<����s�3�|RU��y�W��ϰК��{?|*� ����w��1Y�_ YQ_������4�\V���]�z�k�������Ťܛ
�����˗'>�)`�bL:T@���j�捸���H;�2��{W�crJ����j�9"i#�O��f�o�6�^�N��=#�;�I3d��B�+�H�ڽ�څ�q��u��0Km�r�<�x�M�Ө��b9`O��V�
�E�҂��L&�Y3��I`9PkK~�vy7qp⃩�А��`	�ڈ�ņ6���j�x !P�����e?>ݜ��}A $/nR��d)i~��b���8|o�pws���6j��t�,mӾ�������`����J�To�/�I������XѾ�R[�9��
m�R�2ml���.~���CdD �lf�83P��ų��EG��Mۛ��O��*|���O�B���{�L����l�\�~d�� �튔�d� �xjLEY!u׉�r7y�P]�j#I�45�i�*%�}�*�\�EhsH�_����䱽��
+cM�g�05��Qa�K�0�"��I�N�Z�^��5,�9e��sx &�}«z#�<d�,�zg�S��!�������sT�(�)�����:�T��w؛�5�\׾"iZ�����ZE��JnM[�@��)w��H�l���D�i::���F11�=C���l��{�6�*�`)��/�b�7�v�w3�;��8����Z����Nt�uW
���]a��y�qU;� ��PL�rM&�X�^l���s�5�-�'ؼ���g���~�ds/��rJ�X\��V�y�d!Iv��V�4F�^�0�f����q��kGu$7��D����~L�E�q+7�9�*ӹ�����t�C���� s\��0���O�5��ĵ��sqIqlF�.��zAƠt�v:=��uvz�خ�N��S�.=��3��D�7&��n�
��F�#�~l}�'i
o�B� �+H�L����.�&�5�ٌ���<ԓO_h��e2������F�u���],㪡���y"x����d�\`��/��~�u��&=�I{{!s�	irµy_Ĥ�M�0J�ub����K��E���rf����^DJJJd8%�0�M.���+����fo6�C�z�/!�ܥ�T,$�>pT���s����U��wS0�9��<Ѥ]w��n�a��ߓ���'䰌3[�ܿ~?�;s�V1��C�k�C�S�� ��$)��{6VȝF��n-~!c@��Y�Y���l�櫇�o�/��h6��橩+ �%��4�m�q	1�����|�~l?�n5Oh>�Z��x���՞D���_��[d@����ߔkkl�I~��ϢoW��4���Z&q|`�ϋVnH֖�$����yӄ��c,�û'�T���E��9��U�l�Hy>���F!��X\�C�g�@	��m�҂eI����c�jrʵ��ˮ��Aw {O6��^ql�U��^8s/��-Ȝ�+ȊQ�W
%����	*��=)�����J�B�x��y�հ&��Uӕ�c�_L>��E���^FLg���1I�i��n��G9��؇�g�dX��ԕ1�V3U�яٳ=s�b�c�`֫{�^�NF����KYʨ�ӭ6ey��i�)��=��'kG�����Qn���{����N�r�A(���s�@-ほ�+������[�솝:�d	L�BӜ�9�� ��\G��\9]�g���wn鍏����/�L�>�{�>��|4߫��j�!�,j���c��S%��M/h�}���;�6#��3�zhk�Ws��<UV�m��7�hb�"P�.��E��[��Tf�ӻ�P�<�} �*���MjfxB=���L �l���+�ȈPo�%����_:4����3H0^���c}�ڭal�_�հ��nP�ͼ���.������n�x�
?����/-a�c<���k�ks"uȫ;s�Y����:ȟ��p��Kt�u��>*p#�\�Z�p%_>)Ql����x���#ϳ%�W3��f��_�`�N�)Y{���.�(T��;m76�>�q����3`n=��m�
ڬ���|z���pc�C3�.[�d��I�HW�c�}]Yʑ5�\d(�� ���S�?28'6 ?��e�K�`=`k5�H�{v���f��M&�����ZE�balEaj*3_hX{�V�̌V(q����6n� �2Gv8#�4����W6]���lv�z ��R>N�
�b�ܗ����S��<U��ɻs���1���:ås~z�e�RfIM�cޜ��j��R�\�u�I�rr���,�!�kAP+0b�bι�������y9�R�t59ӏ2fr"(��E�W�tLؘ�쐮��WT-��lu�1U�y�<{��Tf��7���o��� ��������1�YFcƚ��C���r���w[h�X���U��n�n(��'�'�����f5f� U�q.�4{����:z��3��d�}��"�0mzpu�mO(���æDm_D\2 ���;�B� W�H���F.F����;�_\I{)���̪���˼O�]n�b����
H��:E7�˷[�X�# �
P}�N����<{�U�\�s?{y��ؒPC�<��,�&��UJ��@*%�8gv��uc�<�뗄*������a�g�j��\Qٱ��೙�����R�wF�m��40?�Cl))o�����`+6�f�6�L���cP�ic3^���Y|Λv�=��D��]���|&�Z8gc�B��F��s<����P@n
W�x.�hi���U	o3E�H��S	����SuRIA���6�=�΍�Sq����Ԫ�p�c�)���9��Q�Q.!8�]�v@_�refEj�M�3�>���*�6�l�:Ru$�r���*�!�����V��4��[\��ɐ��w�ә�N*����4�IF[���:٩�l^�F3�'�׿��	�*]��zN�ոnS��\�Cբ������:���4e��X���M%Bt����$*��n.���X�K�?��:s&��ӟ��R�K���k�e46A��zė�C#P�gu��j� a��_�����"鑒��(��þ�`��������$��_��Ԉ�7�B��X��w]W6]��e��� ;T$6�q1��l]sjC��&n�u=��צB� ���)�c�����4&��[6�g	ej܁�@ �X�ȘA!h�P|3翍hQ�n�G�xu��@��[��j2{��l9�W�?���P�L{����z�i7���Ź�H��5�
f��&؆��x
Jm��VI�+��N�����Y�����{=�}����Jٶ?�j��r,n�u9ص�#�A� ��2����t|F�T���y-�����V���{��V?+m�4NO�A?h$ L�p��U����>�m�^.�S�"�̇��LvW�Z�c�ֺ���\u�$
��6�%#K�Q dU'(~%���\����'��"��f�T�����O$kL�x�8�AUA0�v��>��u.�Zԇ�~_��D渜�X�쬼�q�]�cLeaGc�L��g�g�!�� u�e[���מ�7{d�nL-7��4�Ue�p����Z8�~�������w�� ���䜭�H���U�S�k5�T}�Vٟ����;P�Gv_�+Xa76�}�A����nD���CU-*�5Z��]"��9❁�/I�<T��>'�
���b�gYq�;��2�W�`9���&��I��C,Hثē~*�J<�JƿD�x��1��Y�{��붧�Θ�TCzu��Oo����ǘ$�j}������V�=; b�"�����kI6�V"��y��*F+������	&�� ��~��b_j�"�k����eʩ��V�ŷL.�\=(PZiHA/��?��s��nO]��R�]�R����B����)�8��;#��/�t���"}3~U��$��KcM�;�r,�Fo��5�-�ˎ:�A���A#� /d		Ji�6(�Б���N
��v��+	����^��S�5!g�VvWV2�)�Y��We`�<������:y��B[2��M����7y�����jV1v~��M^��n�^ �B�g�0�NASc
��Ӓ�M�T�ڲlj�?uڶ�z���hk>.�ڻ#�[ڨ���o�*5X�W_|�g���:u0�?_	é���v�!&"C����{�qx�A�����w'�N�FN
A�����H��#�cktwY�W0`��NBD]���0�8����顃�@�n�&����'��)=�$F�'`�Oӭ�+��ސ��i�P�� �����7�AS��m�n¯��H[������?�>4����Is�h���r�����D)���`{M�5j���N��fG�z�������\��ޅ��z��B4IA����}[�/�����K����6��U�@�f�g�
dN�\N�yߵҶx�o����΋I`��n=��r����6Y��ݱ&��<����R�{�j�
���j�����F "'bq�ރ^�(�-���H+��mS%�*�/D�����2Om�:��l�o ,aj��{�KL�[��+O9�O���'�:�Vo&ݔs2�ͣ����[���=�q �E��d��C�Z��25�k��Ƨ�{�2��� ���aH�/��� u�o�B��3�i~n�Vf+}�?�;��[�@�����ZW���#^���Pzv�>�=:z5_Vy��T�b�	qh�c�(o��.�YOX�b~4����˕��@�0w�&U��%��ά ����qj�ګ��		��q�_'d��ղ���W���p�Ũ��<7׽��>6����?�yS�+�#(��}8��7��(U7Ve�w��d�� L�L_��J������O)��6���#�[ͪ��T��V{���Mп�0��7u\g+f7
퀑��cԘgeӌΓr��F�r�e�?_:�4PE֛FΆ����K{�'���3�����m�P�ϦE�x�*�k�.a��C�Xŵ��� +�j`f�]���%�jp�)�:dc	�@��wЅ^�y������t�_G��g;�[ozj�f��U��_��G<���ϰ_��TA��59�'��� ��KJ�{���G�`��q{+��T��.vw;�ٱ
��3�0�II�HR՛>��S�V%�@�B'w���ȯYBV�g7Q��A8!P�!��q�L�K���Щ9�9m�Ӂ�5��壮��D�7���惒y�d���Զ �6�퍄E��X�J�;ee3�;뼛�S����<�P�?�Ʈ=4ͫZ԰8��N�jN[��J��Gz���o�Ō[����!
aY2�?�TD8���4]1	�����_:C�.��v�kP������K�_�Ģ����tb꣝�zFtS����H��s�җ�*+{����O�a�H��S��:���Nb����I�G��\r~�\٪j���}nW^Ch�M�jif�lɹ1a�p��i=�)^O�����'���.���W�BF� ��vk;:+�b�j׀�`P�E	a�R���Fv\ߺ$�[�|��2����N]y�Sf�rYb��C�[/7�q)������S��_�t�š���nB���lN�9��O�ĩ�~y[P��&������J���^	E������4	����ou�~/�V'����={ߝ݄�h���{��Ģsv�NǴ��$V}�%μ���J7Kw��6��a9`BRO�`��4�E�����瘖?�nOۖ�Y�ӿ��آԘ�$|���
KG��0z����5������N���c�Ϳ,�:����y8��,F-C��ԌT�5��%�������8�3g�`M=�M�G%�qu��!��T�����2uj��܋]j�6X�tb���}��x�c9_��#�FC���y~�_�U÷��te�$����pNi ��'=�m���T����J#����n����_����2�fڋ�;oPL��UmjX�ׄ�'�1җ&���w�ˋX��Іŋ��<��sخ��-�1q0f�:�E��Ǩ�Ldl����щ�1"�n�u�]v��aaU�NCI�?�9-B��S����WS@���3u+��k�L���4�b!���ի�j���S3R
��e�r�?��q �}�	������U�[X��&���BW�ܒ��� ���e��A|i��x`X��O8�Ar�D�T�#�����q4�q�w[��J�o+�x,�m�{����n�%d�Б�����Ā(��]�Z4��W���$�>��RP�K���R��G�z���i�"�Dl^���D¯�n���-5b�^�O�j��K=4�2��R���6�x�SU	C�h��̹ӋVd6�]��}�.��E8m���R&��엽 ����}���"3}�,�$�N��l�{�<�e��|�}X�PbP�/�ӛ�j৆x'��RƇ��U޷ｍ^P�Y��ɿ��uN(�!0�7N,�sF*�e6@�q�o@��÷b�<n�w�tו�Xȋ���d��������-X��R�&^�����iU��_S�p?���#��ј�)�7�%�jg�ɛPo:��e�،zD�@�*r����K����v��+�N=3�x�<� m��g��'Ei|��y1p����u�ݳg-�=K߹������h�X�����VW&�s�DGk�Vι��Ea/�l�V�U%�:��Ja��-@�OD�ϔsħo'���͡��}��gDG |�s�p<I�"�lˍ"V���1��?��G�;t�u��&�a�xao����O/�G�Wr#YP��W���$��|J�F�+�ȥ 5H�n�iE�8)ʬ�*B�I\�v)����K�<����=��jT]�t��X`r�@	d�t�*�j_ xd�DQ�cڛ�q~\3{.eTnl9���/r�p���k!7b�~��Q�#{�Y�5�G��Fߞ=��fK�� `8^p����J�}KYcO?�	��|�;�D����"=���f{�j��.����ט�����=B�P�glun(���S�|��U�YrZ_�j����KbS�o���K�A�R��.�Ɛ<��_�:#�vw��7P�$���O�}<� �7����EzMdBt�`�({u��E�%���}�&&�zV+�)kk�XƍsW#]���2['��aхnŨ���>�%<������Kǩz	��ƶ6�	��!Ju>,�_��;��O$PPup2"C�	:�0�^ ��C�].b���q1Kz�h��l��=S=����}��`�:Lx�����0��P�w8q�y�����%vz��w0��L`)`�~« ]���F@W� ��\$~=|˘�z�"qX̏���An��ű�'M��m��nm�9�y�� ���uR�ܪL��\�i���ߋ�{@��ҭσ�?.2ڣ2�	��C=in���Y��B$�q��1��6�F.�}�X���p�ϐ�~��ۧ[mvP�]�	�����aTG^�K;�c����X�B��`�`���-Ŕ�V8�*H	eC���<f6���F��@܈��wٖ�~q��G����f�4q�kw�������֎G�%O ح�d�Y%x�-�D�Q�|�P��~N����c&Ϻ�XL�����V����ɳ@���fS8�2t�~q������cs�U4��P�U�w��_j ���.C��hD����>\�\�T�Q;�z���npH|ƭ�R�^e�3 |��B�<��>��u�a�B��^ɏ�hv�G�W����n)"�QԮ/��8B-d$�����Fv/4�����J��~��LoCH;V�s����۳��$7Tq����<E�c��-���A;���hY\�)6k��C�� �8ؽ>s|�v�˓o�^�}c���*��ph��Z6c��&�-F�\����eϡC��{�ԑ�p�U@➢J -�o�"/#�)�46���}I�w�5m�,Y�1�����-���� <���v)�*���q�f�@��@z�� �J�ti;7fGȫi�U�xL�a�j*���a�Wa��5�3�5�gT����N�ԲCN~�g���t�c�a��m��]'��[�
:`�#e�
��m*/(kk�����ۑ���د_���y�bGh﹯^�k�y��<�H.�'&b���&W����H7Em�i ?���3�l:)-�Fg��	i��,ɇ!�k8
Ɏ���'�V��TSgg�t�b��]�ܯa�#�h'��z4��~�3K`~u<���"��2fa:6W�����Cl$a<��-!�z��5ם�l�[v{�4��)��������N��~C��
*0���	�g�x�%3�/+�Qf��N��G����PPU��������i�H6Q�����l��%����Y�і}�>o��S�� 91�q�4s�� ���XF���o��MVAq�kʜ@�z�܃ni�r�`�'{�@M@����4vTW{}���6FQ�Sߚ#�~�o
:����X4�e����<�=�G!�ȯ��b�e���HH���m��X�H���K�?���s M~A�����-Ó��@�t��O�0�n���W����ړm�7S��}|*%�W�g����/��G+5���̪���<�S]�7��K���`t�x�����u��|���F�.���&='߱�>�gO���!x'�`���g�/d4�:�����]�b��%�:&���#�;<	:��}ۑ��x�+"IL�����5�ǀD���^�,J;j=�nr�)��?v��Z�t��1��a�?��K�b�c��*�(�l�������v�6������{�`"b�ƌ( ��My�~�gh׼�i���%]�<��ڒ���it��_	G����_)�M5�
���JYɱ� "�շ_;1�U S�5�3�PzU��K��:��(����ͣ�(̻芩�'NiPg�s?^�I�`�MIá"���8|q��Ô�P� ��b�Ǚ��aY�"Y]�:�ٖ����a��}�y{T��S��1��L �]
�,���9Z;
m��ĺ��� T �4���֭_zD�L��(��K�D�q�G�?l��А�?���P\.T�U1E���l5�`��+�n�<�UfR�~�B'�g�9�Pci�E�/�Q�[��r���3�?���︌�����V�=�61��U�A{� h8O�?k�aZ�/�g�2�C��4k="Q���e���R�BG��Vk�x�D����}��%A���+�_��X��;��Ӽ<�ao%�i&v��T1w1��c�	�S=�:�����Q}�>����P�O���C��~.�R�t�6=�&{���^.o��z���G�@;�.d���z��xh��
�_��E@I�ɴӠN����حpm�n�*DP��'"9���Ϲ�~)���X	�	�7c/x�?.���Z9;p�Y't���i�֦��e�ũ>Q�DI7�AL�l,1vy+���U�K<e���i���6m�G�J~�ި��i̪7�>u� ��>'m�8,���k�]D�m�n׺UY���ÉӃ�޾�{9�����us��c�)�ͨт_�D�܎lʉ=��}�at~bf&��DM� L� Ŀ������s��������K����zn};�y�^��p^���D8}�ت:��� ��jⲥf�<�Y ��&�q���O�n�4�\:qɳ�����;�!��L]=n�޾O�A����]Z�®��u�����b=��4�ßSi����!�x/�`|d"��������ƌc�W�Sı䶠�����Ƴ`�9�Ӻ��i�s�S��`�+�¤z�8BGQ-����DzxX%ou��fR��G�dKeWa��������������!�I�XN����8|/p3f@#��' ��
C���n��7\L�i>�(g�M��IE58�ܭ
�:ni^^�w��E�_�}�ݛ������ȝ�h�n��2c3J��G�}�(E�e5EF��ـT�9���V3��������)X]�7Bb�u�3�⹧�$���C��� 0<����I/�~8=[vz4LE�^mpt|��z/����<�I��;���̩�wӱl���@�U�zߠ�����dP��bDM:G�H��V�2\`�٢+W7J0���R��-��.�*�����e��AFO�PP�ꌮȾ��J8���2�G_Ei�,���?ܽ{��TI�c8�+3\JZ���d�u)����Gh<i����P�G��7�ި�����ZG��>�O��C?�L�1�#�t }�r}�>�hC,/n��b��<�Y�����Q�I l�mU��ſvy��x��خ ��Vz-�/0x,���Vg�4�j|�]�r��������q�,=�#��m���i��(��.K�X���/!���l�n���~��3�p�Yo�G�����jk �IBٸGN���9��8~&�����_���y�C�ToX�,p�l%!�� ��r��C��מSi������)�=�3U����'�W����������"����Q���ܥ��D	(�n����1G��̀T����p����0��Mfx?O\�� ��K&�b��{*W��f�oD�3�܇��Z9<Y�9N�P�f{�XF���� ��W�����d/*�CْvMMA��ܽPO�������?^&^���C���m�o��T�9�N<��G����s�է���������'��z���ٷ��XF���SP���&�<��a�@œ���I&�&PQ���$-�]'#q,Q�N��A'��#�򊋽�'^��g*���n�r�K�H<'`x��j��r(�ˮ:Z����P'
A!@�~ߡ~^���s�����d��sxa��8����8�{r�Y�g�n��#w�R��+�U`�4�0���_�E���l�2g݇:r�u�_�$e��4�Ī���E��������H�Y1[ޚ�����<��y����i�/�y�(5���Y�D�Ϭ�z�1���j�P�	G��X6�o+�=��#���e�|�Ъ��R!���r���,�Tǌ�#"�?d2h�ٟ-n����1A~>u���u��z,hEAb�3�T~����T�U�Pp<o��oI`�<{�E�9�Ӫ������0U��D��c����r���n���K�B)h�tr/���Ka��G��h��xX�o[�,>�>�z0�?�����FC���T�뜪g�8yߩ��*n0�7A:��oZ:=�i�}쿉�"4n#Ԣ�r�%����bE��=�O�u'�D�? ��N�==�a�ݵvV�]T�)���
Q}h��M��֏�i�J�^sH`e鍽�]���ˁ�qeC���&0�2����.d��R#错b�t������xM��Ǌ\���b^�����_W�?[��j�sn4w�#3��;����9�1 �}8�4�.g�L�'����8���6^J����W����~ח�Dm���:k�}E��r�=i�w��ꗦ�F��:�ʞd�T	�.Z���{�u/�2���s�Xs�X�ԕ�9�����D�K5C�8����u�u�V$��ko���7�r��yv>��':̼P6M��x�x.�K�0�Ƀ�W.'�Ϋ������&��ۖc�S�6��T�ODY�ž�Cݶ�M�h��;�J*1z��P׊W�?�k[��	��}��[����|q�9��R|Э�4�r��)f<�eH��ӥ�Vƥv+��>�H��c�i/���F���ng6���`x�t0}�a��H)���ڣ�b�R���9h�B���U��}���ߛ�����+��:��m^��e��[n�(���u����ߜ���')ٺW�ڦ�E���@|l�^�J��<ڏa��O=a?K��ti���g:1ׁ��`�8�'��{�b�qy��T�^��:��ؕ7���<�3���a�&�w6�Uk�oO��n�M��������V�q�_9�$��@bd�l���~�{o4�G�]S͑՜9����C��γnQ;?�3Ψ�b0:���j=>go���J�ԩ�y ������Ȼ`�L_X�$��=/8�ỵ�'�7p]��OK����U2͑����q�`zL�ã{�[�U����� "ǉ��w����%��ը�ٰ0��H(���}�g��R�_�o�:�K�p��X�j���
�-� ?��"4�skS$P�����������?�Tθ�"��|��t(�h����首��J L�K|�}��1I9��T���!-��B�&ibb׻2t��ֺ��Ɛ�a��Ҵ�d�2&m�&J#kC>H+��]����>�N���a�B�%X]l#F/��j.}�17�C$e'��E}c Xo]�������QK]!�E�0���Q�unk*!Z��#2yK�� �ź��;ɋ�f�c��-�j%-��iZ��
�Ȣ�ǽS]-@���^�b=�@�j�?,�����`��Y#�h@��G�ygښZ���?
��In�a��+r��Eb��w�x�I9��s��8r�w!�ȰX}"�{��B��gْK�H��|x��m�F�X̊��3��:[-�d#ơ��:;m�H����3j9h؆6B�����E��צi*. ̟ս��E�8_nִ߳X[Xgbx����-I����c��czlupSi�L�����ZjsM�UR:�4��Q�_�}<��z|�M�9Xd"����U��);�=�y���uK� �;��`0�7�V��]I��� H�,g$AFL�r�ޏT�"�+΀{i�����
���.��6\'숥����sw�2r���4K�ۦ��\J �V7?��<��[��w'�
��3����H�$����g�\�?�  x����t�J-~�f���M~���b��\���Ŗ<VN䤩:�jy��&7�f���P��g6b7�m�r�b��^=�Eh�_P*Ԛ����������ح���{A�W�;k�9 ؽ�1��	�ټ��"��?+�~NG�y�.p-&`��8�� $�7��7�*�ZU�����[,)��w�F�&����D��	i�Lt���(�%����� ��ɋω\�_w+���xg�aĮ����l�1Ƙ��\+a,%tR����;B�;[zEǇ0/N�����P\N��i�P�G�y���Mm��Z��[L��i�ÙP���wZj����Ȑ@R����y%���sA(��'�\���̥�4E����U�ZW�'k���[|ν	���T��y�����Jg�����n��-�[E!n�z�zKGu�r�wLy���b4��(<����K^g�]G��)Lq������W�Kso�E�.g&rK�5T��������:�SRRAk�hG�?eT�w%�h�+L�_�����ۙ!>�嵚�z]��&Xo���讐Jc��\��`��ڵ)`�X[Th[ѹ��B�J�Z�*���T��tl��>{�Ჟ����-�H�KF)[h�;ܦ��1_X6�W/R�\��\�
%��ώK�r��L��"������vr�K��d�&�`o�������=�4g� �f�s��&<�Z��Ǎ���U8�6A5�r_�������_���.�3���cDʵ�Ō� "^N eK��f��ܔ��~���tk��������W����0�4wu=HI�л3���x������#��`C��i6��}UP׸�hV��)]_�������[��Wt�#����x���f��	}�'��b���N��/�b\�a8�G��~�w���p�U�\2f�׾�g��<����7k���c���^�2h�>�B�Q�*��ƭ��/�[�L5���?u�fi>����B�\��Ҋl���e$:87�!l�T���߰.���<�p~
�t�I��������sہ[Jr�V� x�f-6x%�p=��uxή9;���3�k��o�C��nሜ�5�2����%l�Ur����9*Fi� e gW���#��j�H3������q�w�i�O����_�w�u%BE�9���DiW ��D�)�ǧhj��a�#Y
;��%s���^�O	���V%Z�Oe�gU�=�<tn�?�������˯z4�Tn�C��ɡ��Z���1y4�o�[L�H�p��}]��4K3�p� ���r�g3�6
V��ч=2�h� �?�.Ֆ����"´�gV��"SL狼�+kk����4w&������%jo� ��pӸ���^�C`%g^"[?qT�A(HD{�|o4��e`�u˺u�{kS&le�l@� M�M��G�<$&'_͊F�	��U��~Z�
-����e-��j��tx��hi_f��H���AGN�e��Rϸ������Ts�~w$\�� ����Z`����s�tn(�#��� (F�OdQiή�3�\kt��<��̱T��M����&�ô���C�j?Q�?Z��;t_뒕�G��ࠇ`��~ �AOs�Gj4��9����	L���N����X��G�T��D��D+�u�_Hd��������.clI�3�(Z���%��.x�	��j,@&�M��,�:�Yo�;%��?hO�=Υܜ��@�)ˇ�!���.�ɵJM���b�.>�sX�L���	�����]��^ɑ�?\}���5s����s����<���m[�z�I��cW��NKxAS��N�y�f�}��⸨��Km-��5�
�{�bJ�3{��
&�'���?E"��)X�s@�D�cD�U�P������lvV���a��]���g�\S��E�`�~����P_e�x���δ��y��<+5�A��g�K�,5��^VͲ�l���]2�L@�:K~!`�����I+�~�� GI�%'H$lyk��u�E&���D�^?k��'��a�����y���ʿ�6B�#wf��G����,�zi=�AM�8,K=3}�L���=)��`?����m�'!Ht��9���m�&ȍ�ht.���g(�ʞ�(��^ټ���S5p�]��ZG�\�N�!7� >�Cf�g��<��+�ʷ�)�?8��i���p�kC�Q�)MSZ=����`��	6z�{�0�Q�y�K<@20~�������������V����t�����3gZnq��I��Al=�7#�|L;YZ:��}��n����"{�c�u,�8]!
݄�QŘ�Y=܏f�D<��!'�*o��y�]/���*���,lKd	�C sV2õʮ������L4ە+.r�����)L|=��-��M���Xh
��պ G�k:�}e��<�|Ұկ�1bA[(�9��4K��i���Ol�g�_��I	����&f`>��96�^�����9�cF������c��w�֕5!m?-Q���m�"�ZՋǿ�Dw�u�IH����^�}�՘��K?�@��e�0Xg�s��H�&���O]~�����C�t���o�&�o��!�i�|:}�"[�d�F\���Q���"}��o_i��e�Zv���x'74�W�]�~g��&$^9�ڇ�[6a�_���J���H���}c���j+ל�ZYo�V8I�e��g�}��SůFn��ߖ�"�e� ��Ng�'��T��úW� ��|�/�.&�?���5�h�g*�?E�x���P��������W��-�>��(:�����"�Zz�h���.�S���[8`�yz�L�+�4��>\��U���h}$�5��a�����+����� oNz�in�����l�4����%D/b!FWVЌ���je{M�����O�<R!_[P�^�ہ�9}�Д �E� ۿ��$��y|��9'L$���_Y�3V�����t\��޿C������z0T�Kڪ�M�����0х~k�H��#�C+��RW�FSo�w�(�WM�54q��P �'�lGD�Z -��e��FP\9�]{�������Ϡ����Vƫ����UT�6�L��q�	��&d�X��	���";��>�iw���y����p�q��Ahx� n��wɚP���Yt�m�|
�G#=�y�W!`j�;�u����C5���iD�����6g�tu�&��"d�7�\3���"��z�	� " Nɇ�P��4��R� �&E�{K�H��4(���u�t>1��*w����<E{r̻�j�Y���iq��w��E��yɮ�7{�p ���I��*5��MOG��7�a0G��?:�ݥ��F�A�
 I ?勷�V ��~m�6ȥbh����V�Д=���c@�y�i�X��������Rӥ��}��-�F!��c��ыR 4���e��u�믋0ɿ��zP6�d����}�&�ul���!��ٖU��������5�L�a:�e���+��C�psGV��j����� �*%׊'��2����t�f�[å�M��_ 
[k7�*��0�ȹb���[�](UZ�c��Z1���C��Sp��`��;�޷�0c��o�"��ϺU���ח"���:�+~�����H��`��m�9������u���⪷֤WʹŊٮ�&�0�J0����|�ù���[Y2��;���Os��#����쪴�M������I�ѽ�-�� �0�L���g�n��������b��{	�t�ţ���C�F����I�q�x6���R�j�f�	��x���>X��u{�Cթ��qj�7�VD$���2ʎ^@	���Oj�A镾Ktq���Y^"�w {4��Z�{�)�c�k3�~�����ֵ-�䩔@��+�"���_�~���a��#ڋ�T���g�xRV��.+��׹hc40_�b��G5����`9B�.�I�kׅ
Y����;����灝���U��c�|W5����v����1�D\��4m�.�R��������z�L�t�@�re$gWC���5>�����Aj����p@�P�� 5��3�m���� �Z;hob�����T�?_ �3�0��e����Y�nɳ�i�FO��L���^F`:[�Г���'�
0(��!�``fי)��=�2*!��9��v�K��/v��<1��78\�w�8�?a��:�|�?�ѱNo�>CjDA%��b�+�1������
O�ݪ1��v[`s�����f�c!%�̾��P'���}K�+��-a�bX�I�䆳����cM�|��(6�l���BP&��󕉹s�%�i��k[��J?]�v�+c�R� n�~� ��[�F֚Uo�B����>@��Kej�� ^:c�gi��	r'>�����L��A@t]�3,ƈ��eAJ>�Ek�CZl�!x������\=����W���~����q�ǹD*�YZ˄@�I#@��^w�7cߐU|�V��,jI���]O��2�^y��9�v��z�y�;�Tw}���co(��5n�OwW���lF��'P����lEV��Z����iI�>�C��ճB�{{4�Q�7��2��԰L5w�4f-q µK�,<E#��xB���wb��Ʉ��}�Oz~������f�šN"���3���0^�R�6J�a�w�тu�t�.��;��.����aR����y:�p�*�n��B��vۅ�����#uga0������ήÍz��N �ډE,|�Zp_��1�ɐh)�(�[BYW*��p�"PK&��(`I��څ�}�x�lzɨ�e����+������Y	J�ox��ЬP���<S�e�ф,��4{��t��m���Z���r��9�\P��S`��F��ߓ$��pso�;h��(���M����<\eXT]D@���C��C�N鮡CQAR:�����:���|���<23��Zk��F��.���m��öNꮨ��j��XT�j��5,���x��.���L�,Z<�eG��oQM�,�������B�_��On�1���$"ҤX�� ]���x�6����@��g�� �s����
���(u�a$���O�&�9��݁���ql6�C�����P)���n}8����qU?ȕ��`��f�㨷r���5��p�<:�ڍ�9�@�Ӧ^KY�4c�;!&�Gv�@�[�p.B�aN�Cy��-�ʥ}�Y2����c�W�(ZS&���������=�@�#�3��R~������WA@�,�,�h$F��P���J �_���8�ʡ4)ܑ�������UE��ʡt����������P�Ii��5_�;x���hc��)?��|8��F��]�~��5�K<f�� �J���F�]݄ÿºiD��V ��ih���DĜ�� +N�H��,��i,p�}N!¬������P�
-�D®���%�жj�.�54X�h9�@ ��k�փ��Xy�P�2@ުr˘=�� ^��"�T��[�tfh��ه�G��Z������]a����ԟ� e��qڕ�{�������5w�Pn%B`Y0p�;�T־6\��
��U�L�&�� �t� ЄWi�QaΓ@X]n�S�]��'o%����oM��3��s�ZI���`h3g��Y�;=����K�?t��n��U&�Ո(��xx�Uc��" ��E�\.�vZq�ȗ��#�n�%:��
l�@���`��Py��鳅�X~��ž��3r ��b«x6!&Q���
� ��g{�΄7�wt���b�H~����i+�3%�Q;��X���sz�S<E �w+�_f�py���@aK=$� ��5j��J��	���a�V�2����|�a�X��Jzu��X9�}i�V�M��v�g2�K��p�S�^�ҜN�i7��d����;y_n^�����!������!3�� ��x, -�(�G>�	?���~ǚ�78:! �\���0�8c����w��]�P���^E;�E�$�+&G`XT�^L��![1
�!���C�M h�t�;v#�~S��@ .��I`��#%�=`��i����Dɝ4�>�rΕ�.>�Gb�]��óNw�r<�4Ϝ�2�������������6-�T�����S=����	��C%��OkD�}-j�`�5г�a�̌�<-:��g��B��8ؐ���r0*�^�Ċ~�QȀ��_��v��:i��\������������99Z���t���s�4���iK����hxI�S[-K��$�
��R�����/�V#}�d��Ԟ�v�wsv�3[���Co��˺m:�S����~Q�+���[����unU.�@NP����JM��ͮ@;�J��}�����=a��&��f�3��9bv���m� ��L>/��swS�'�c7���G�f����&F�%Lu����v8�A��CYK{�I��g��F3�� 	"�u������x�� $�G�z>Z��ɰ��jA�6J �ӱ�d|�<�Z��c	�������'����2��:(}3ш4���CP��62A3���E�-��q�3��d>QXVh@�@��F�K�o��?N�M�YPpe0	`����h0�߰0:�Q�^�O>�h�&a��Q,e�.�4���O�Y�*�f�J����PRp���N����P�L�Y�$B��y5�%ܓf�i���=��?^�ץ%ǎfR�6���j�
X׈�U}��u�+>M������l�L-|o�	l�����g�I~��6	�ƺ�5˪3�������ԀH0������w�*�,�a�C/�+�w�� Q�U-��w����p��Ӡ���t�%r�n�=��uI��r��ڇ���D �h����+����A{-�~��U %��T��hB�S��!�|��"�gm�azy)4ɞ��*�f�ƽ ��r�.�0�pe+8����b��zu�z:x�b��{u��r[��jk�oe� ���_U�b^�d%����61��7b05�1N�g�������S�J�v� ����g�=*6h-!���������'�.�l?�����?���N!
iue��po�w2Y�>���a[^�hT�d&sR��lB�ȧ� ��'��Q�c�S �����#
Ni��#:�l����\�}'y�d� )\�����ݤ,t���2��1�^���)A.l��
���UR���(8������b��zqV��I)�8И�'����u�f#���p(��S]���hI��kE ��u� �=-^Xb�EQ&\ɂ�9
�� ��q���PQ����eHJ��q�>dJQ�Ӂ�+,�z�8Dt�/�d cX�Ͳ�x�5���q����?跴��zJ��m ��]�*8t�`}�JsS�W�ju�q�<��$.{~��o����w�?�G@`q~�;�{�:,�h���^�-C��b�B�< M���h��Ø��O�O'�>�zQO
�|�"#K5��1E�C��*��ů�f��q�Ѿ3a;zG���yDwБi]/�V�ڭ�\�����~?��K}���� ���E�|7�hH/�8���.����]��;뫦�`s�V4�]EA��hHzx#��&��`�����D�ܜ
,U��W:8�{�]���38�TU�d>>�y��b�$(</a��-'��(YOXl<�_}}�q���5�T|����ER�l��r㩹7��3�D���i����d"͈ՙ&�^v����g�Dw})��g e.���d��x�\0{��v�xZ� �OL�uF�H��0y�\��l�Ȃv�����V�p7T�� [���5{�t���"Y�M3�>
~����|x�^P����3�'{(����^��8�<�2EU͡�)����� �|(|���n��0М��U�{��.��+��A"
i�G�B-ஒ��8��p��7�jm���?�Ϲ�����[�ħsa��+}���
�-/�V��c�L����`qu�C~7�*0�$��.@��7f�?�O�n�����Y���:�[���X���������s�[@؇����	��C���o$���N�-V [pd<���}�[�x3��>M߻��dQ�K���0�.�b_�~�2�"����F���}gތʽ/�H��v=���l���� {� P/Uiף �����	P��ۏ��.�8��E����]Y��h+q���w��/#�����?@������������mMBy��Z�����F��K=�q4��^=� ,)� _V���?��;z�Ԥ�?QsZ�00~��
�咼��?k 2�A���$�{���~���l���[�
)�c�?��{��6��kh��K\�0� �4�����&Μ|��+�����J��J����P�#��u����L<��<P��x��(l��wi1嬜-�)i�A����v��V����h��˭�*xl=S�;Ҏ��cUmt�W��JU���[� ������!Q���v��e�iS�e��zpLl�j��¬4.>���=���hO�-t1�j���;^H-}(����k2&{���������P++r'e�F=��8*���w�6�F�N5�m�V�_�ُS�\�ϛ��r�z������$x��ċwmK��[�p��L����ݻ�]�s��C�a��iSZ}�E�O+:oz6��9�&H5{oX
p�����/��5v"x��>�e`��7SSt��(�o1�ї3�n[]�D����*���H~��ϲ��ϧ�� |U�!�%�ǡYۍ.���yn�Lw����xe~Uw�G�e'��˩�H����f��Q8^��"c&c�gyΛ���c�hgY�i���!�3Y �n��~E��$�06��0[�"����E �1���ڪ+�xO�p�%����M^qކ%�)\��w<J\�n�w���	�W��)5ԗ����K�2�B̎ ��P+ߦdV�'��}/⋻�P�)���ZJ��C����aSՖ}c�l�O�ǨZKɷ��jrfS���<~���}/���ϑ�uQ�>*��ΟH��5d����bRR�,RR8kUۘS?za��L�8�h�
N��w}z55�Ng��d/��\�@f�ШITe�P������n��Ȼ)� 9�of��X>��E�؞:Z����<*]�~s}�|7W�j��	��zV�6�> $Z��[薋~(�p�i�U���l����=}��D��;�<t�A�\�VY�Ӳ�7f���!��>�Eh��NKW{J�������gf??����FŞ\��W��ۓt��<б�
�8��>Q�V��	VE�fzE��!������$8׭o,�jX>p�X/ѲC%�J�����U�*�2I���	�]7��?�|twG �ج�z_9�ǎg2fY]��t�r��1����L��k�=�d&�u�P��\�J���y]����q����(���tw���V~�W���f�#i��Tpdd.�����om��M�����4��
��6z�J�0u\<t��O��lmK<c�߭�����(��q�P\	�g+W��"�P���X����#1��)��x2>Ńm�9�ĭH?s"��a(�LF��~���y?vf@4��un����1Y�x}*S��L�''�����!����A�
�F�V;߯��G@����b���� v��^�C�Z��nB�-&��>�H3��P)u	�����a��s�RK��t�	Rms=ˮZ"
��?���jjs���5�I�a���F���q���d�A~��� �N���giQ[������;v�S'��or���U�A8Ɍ�-�=�X���?Z(�x�%i-*���y!� y,[q6)��X"=����X���q8v�<Z݊���/��y������	%�>3���Q��+�n���%�C����w�]b�����+$j�����r�uu�
EQ+��5��F�qَԽ��1�>����E�_ib�k:魏���_�@�t�/~e(k!�{G��ä���iP�WVWI���y���G/��ٝ�v7F�T�=��UM�%AhJ͂���s�W���>!�T�L������HN
���w{��9ك��NHM��>R�9*�o>�i!m6�k��>����>���j�(��v���W�s�L�A��AM~�/����W�r3�يi���r��#�̢xS�WF ����8b-����u<͕��<P���Q�Sٺx[k���8MI���i�j��?�Uq��Gl�s0,�ʺw�GF^��J���A�hs�FSP�8@��\ǭؚ��k��&	D	��W�f�g��9*x�����f<���8��fc�N���ji1������O|�s�滹���q2���N�"����\�zJd���dD�* .5���,V@�.���?����2�\H�\����SRT'=�啕�^6�ϗ7l��!���9TV?r��&[��Gw���u�g���V�}�,L�^/=�jفv^�Щ%x��d�m���D��̭��ܾYVV�����Z M�5M?��^u�6�����~�Y�*��5d�HF#�\�>>���V��L#��4w�lIP�{��v�	���� 	��W":?�D$l���w�a2��sTO��X�f\Чz�tA���^#���-͂�Fr��s�[��%o�`4`e3����Y��J��,��z���t��02*�}���qt�{�Hg����q�o�]y�É��P����]W��ĴZ�c����nGf�<���}���H�_#bw�(M]/�yr�d��I�U��l�sx����tnH�۴m���ї�!9=y�;��s�������a��R�Ob�Aq��Y5>�y;��VnX�����6�$al����&�x�r)&�0蠥�V���SԞ]�B��ʼ���ԶU��|,��E�$��c��KV,b}1�c�$i�[�zQa�<���Ȯ���~��GI=�n�HӲ3O�K�����p����dio
��4�Lu�F����������]���9ţ.�� �P�I =�"�,��l�z�,�v���a%��43oe@$<C��-�V�3%�����%�Ʋ���֤��Ws5����;�W�y����|�u�8әܻ�ժ�E ��Nkd�j�nƖC{5���wM��`V�H+aF�п�y�vva�GKC%��ﯼ�a����T�KA�)�pF�� snC�*�6�hr��K�����9Q���(�1��,2+iH���
��͒��9u�FѠCr[����it���B
<,۪�RpJZ�W�)�n����c���K64��f!%��o�2>�`���h&f�7cG���N�w)T�{�M0,� "DENw�s��l���߮@�Ϻ�+5S��d%�I��>5L�w\3��F��]�RX�$ƭ�l���P�tLgM}$�Jz����M��"��TGB�6cpP�d�ShEq��.�����
�B��Z��gtnkc���Y-U�����n�*���o��_��U�I�x�H  ^�J7T�Si�k�۪����ZΗ��ŧ�!��9����k-�v�t*��=�!!Q����9|%���C� "����B�K���6��-��5���������bn��7�9�'?t�<Jt����\SD}�iV�48�vZ�F_��WM'ڮ���8�3��p-c�)�-��D�X���L+/t�}��['s5�qy7ݷ_�ĝ��ʌ/�JV��U܉�ۋ�E�{�|�9�`�pbb')�3sL��Ƭ����@,{������_j����(��:F���g���7
�@+���y
�`4�e
}�r���k�)�e����f($��oBf<h���ڪ�곅�\YZ+�}f-ڔ��w�C��i��N�W��W�v��Xw�q�à�XOz������1##�����,}���@����~��6��ʙ�;���.��?�MZ�7A�	�T��H������X�5�U������?������44ߨ����\UD]�г�UIB��֟[��!��y��*���]�q��nG�s�32�C��C�����ed$���K�8W�W��㎵k�^��j�ɭ��	��ThD�e��[�ݎ��^�)�����~�{;bl&7k�߉RT>��pR��(֎�z�m �;�[�+�\�4D���Q�0m4ꃏs��,�Q�R�-���}��n���g�����؄w�=���d���E�7[���?�k�_���A�4~��Ay��">��Jܰ�v��]�[i�j͚�`�C��[��|墘�bMO�ϥ"5�_,�ln��������u��RI�0��^Z��;C�y{����7��ƌ�<���!���W���VG��[I��C���/M@�AKG�_%Ռ����w�F�͔���/�tPFg��|�͓/f�>�̷Y�i�i�e
��K�-��L�(E�����y7E�s�~@���������p�P-�pyW����]�+
5i���e�Fo{7����0�LO���C���=���/N�4�j���o����@z���˳��̲���jKB��3-*e���T Ŏ��Y�:g��;�VG9DS(����$c^g��Lߦ�#�3d��%{�F����*��#"l����D�����s�g�J�Y꾧��l�ˀ�{R��Ҏ<��sC�K��(����[Y���2���O+��V(����ɻ��Z��� Y���g%6�\�y��hZ.6�y~����xGU�W˪���js�3�׼���A]�>���p�p�N���Ե^��"�;Ȁ�/��.` ./@K���,�}��=��k뢝w�����!���\ܞz�&Ü�.��ee�O(Vsg���e�7�_8��T�����Y����bl��b,70Gs��(�~�ǜ���j�+��e]��H3"��=՝av�܅iT2�ǈ���f���b�djR�/v��ǭ����v1B��U��jm���\mW����Օ� 4tv@�`��Z�i��c�j{G�΁S���pFƸ�op�z��1I/QYmҮD���Y�T�Q��c�����v��������B��;�0��jsc���(h[䜙�r��
���$����Ò����5��)�'����]s3�����
5[4�����A���Կ���:�O�H�F-�a�DV'Y��
,M��2���4��*7�Ѿ�村�{P���S?n�Mq"n;YFB$e[ꡂ��!�͑M���E�{h�̬k}�c��n?���e
�9��h�_�p5JY�
������j�U��<8�-p^�no�̹5E�T�r�<�3�>]cg�2k�*�JuY&������O{nD��Kq?b���3-	=l�7,����(e?:��;x��nL�pQ��W���o�p����,�R����5�F�8M�4܂��	��A��U��ՄJ�ѽ�n!,�I��Lm�i]	�\����������&t�e?�r���KMP�ʳ�J�ѲW�o�d�L0��yD������0z��m�����*�)�&=��,#�*�T��~uŪ;8ay/�MF�Ⳡ��#p�;��ʥ-��V~u�\�ի4ř�|c�/2�1��̫�|�UL��n����P����i-��s��Q�}����݈[#xaf�j��6��aI�'Ǭ���Z���hwp�Lnoo��W��h�֏��Ip�OP�U�m�h��i�8��īs���R��������s���d�m�c����t{�;�z�A�:�~(�/���P���|I�*�c�'}ZS��N��F�N�z#�v��ɺ�[�D���[j?���~uM�地o�w]��HIuE�幫6Pןˍ����Xz
syg��x��F�D-r�r�r[䙙�-�G�
H�z=X����;[o�ڬ���֨��6C��[��BŌ��対�_�lK���F/0��VD�R�lq�~�a���X������G�栧FL��yx��HFG�
ň[�ʇ�q��TQCx��W��┨���12��tW|.�PT��?���p|����G��8j�;	�������TiۙG_�s_�u�&Dcmw�fp�|f�c��6�'���Xo�)FEE�IEPpی����0a�u�AM���:3*�
y0�Ø�ᩣ�0>D�9�|�U�������⭟':`?��P3"�u�8E���[�����ߎ���˕_
+8i_�EUX�c�}uNk�:3D�<{6���jB�ִ�TcU���>7���4���/�
�b�Ep��qثdw��!���~DG��M�&�SnT�T���9�������I�Wr���K՗��x)�}XG�Z)�WjJ��;�n�{�z�p�`n���Fj�{�ݳ/�+����5ii$��8n��x3�}D�sDV�.��;�r�l��M��QN~kC=D-���ه�cx}���l���q\#i4s������&�1�B׋KUȂo���A�_*�����1�2��˯�߮��Ti����yR�����e�ffy泵�崴&���婗�"����v�}j��믬d{a�[.��צ`7�Eb5��d+ڷNMv�PQ{(T{��o��ռ�G$�ITR��=�b��.*���Y)�7���S�q�Gf�"#J�����ѐĲP���#<��~�/�K:��/��=��]���%s,�)�e��\�D�����m�
w!9�@��Ӿt_K���s8�q�*��#wN�)~⑗w����4l$�/7�b�S]\m��nY������y�B&��Po���,�����jP��`�����K��c�-�G	w�&�;�g�)�TCf4��=��^O�45L\�V�����Zn�#w����!	ĬFu:�"-�HSh�`��3 ����;����ZW^Ub��y�=�u��a�k���7p�����?��W�E���h��{A�����M(�r��6�^j��sOn$��n
;wJ��g�$$��|�gN��w3|� 1ЙH=0�ᩜm����'1�wNo"�V��5����ō��e���B���Wz�"�'�ѹė�Q��ѝ�ոR�s�l��ֹ��kWD�NQ߽n��-�s*p������z�y7�hw*�Atb	G�����X��Լ��R��Oj�'�v*npO�V|t5)�����Tu-}hߋ�%t:��h{��qM��G���������K,����B��\���ќ��
��Zd<�36ϗם��.�=f��+�~W2g� 鼓�9��a�t�m�J�t��Ŷ'xD<+)�n6�SBc��!BEW�)I��n���=�Q-	O��}b�(IG�m*(�VT�y�����A�vM<�:�]r��ǈT9����?Od��"��8��
k7���ɓ�Dy���5.cn�)����G;'�/�t����\62/>~��J�'��%�Ԓ����RP����)_�4��6	������ �:>��b��:Zuu�����Z~h/��mg+g��[����\%m)�+"l��8Li�*�MS�{ʞ���D�v��}�O�����	�!\^ݝ������ ����3�����}����?�+9���{d<��O��c��q��D� ��Bhs7|=.)����f�e��r96�A#���O�N��_�u�B9|��~�!�ֹ�T�3�b�g9�(��_"΋�e��8�ً}�]��w<��q�s1��-�G�g��[c��;L��XA��6�q���|w������k)��5)��Rk��X�w����`'�Ks�dv�X2����;o� }Ҧy�v�\��Z����xN��uJ���.���2e)��e;���7��T�0<��s�u�!ꈃ�HƢ�+�[w/�E���ܕ�4H�sn�)��f�qi��B��Գ��d��!�@�n�tWe"��+Gl���e�A��1�8�実O��#��`���2��U]vK���G�� �G�h`@;&{`3����Q���Lf>2~ei-Go�G�o5�fت
Xx�Y*�V�k��!���a/q����Gs�r��3,�nT���uxߛ�w�f8��!;I~�{?r�ǆ�2�����.���)�T5"�Nh[M�%�1!��`��*;6��e��_朴��S����ܟ�8xی)I	���]��G����i��-{�bMJM��/�ǔL��uT��k�;&�����V�͹��m�Y���@��HvsFÁ�iΥ>���$��8����Z/t�)a��B�������YX���ERk��40�}�-�[!�!8l'��shJtz&��m`�MiA�PmE�juJz�c#a��Xr{�D����4f�nI�˫�C�p�����N.'��5Q��>{����p����$�H��Uc���� ل�m�=�\�j���������h�iW�}dDP�^���@(��[y\>]?�>+����l �=�A416�����K 'J��A,�S}̑���ӆa��+���<W%��.y�b��CZqGٕ܏��7뺐i���K���OU�����)o�\� �����GI�r�(�ö��y����d��'�п���+�4=����O�	s4X���W.7���?�z��O���KQ�ud�����2;-�%>6oג���=E[s� p�#��
/�d��6R�'�j@��%M`�&��C�,V���g��j�K�u���n�����s��
�c���v���J�d�O�h�NT���n{�Sf�;��xd47��E�dm��[tK��}����p,�k�$���8�:vDc�z��s|xI��/�3랬2���O���o#�s�uW�L��0yp:>��'lJk&X�2�`�z�5n�Ѐ^��+�G�(J�^v��-v��@���z��]�V奷���e�4���.����nbqƯ��J%�;~��܎*6������k[V�����Ŧ_ ��y�B
�v���K���)���Y�Pyp��U(�{N��X���Z��8{�h�!j^.�9gB����x>���,!.=K0ٻe�BD��bߓr_����
Gf�x������2�(D-�Vu�PF�qi��{�#����E�x�#���,�)o�+G�������=�n?;�!�/�(U�t����a��y�Lpj���Mr����9v�НLD�ˀ<s-�� h�y}ڽ5ö���&<�/u�9}�h�rw:����7,\�h��]/|�lQ�p���c���E,��_TO�����9�G}�z@J̚5�僡C�%A�WC��Kn�����&�e�oMJş��J*r˓.ɱ3ub�d����LT��=��1>��?� 8��~�FS� ��8+P��M��G�� ���� ��|���e�q�� Ũ�[Y�}�W��k�r��C�(-LpԾM��fӨ��.0Zb�W�?�#�-�~��!@��~P*�jT����[�P��Y��X��2�:A2�Kj?�%����`�G7�՚�gߚiA�s��ZZA�w��ȿrW{�{b��.5R���x�%@��=�޽��
T�(Ʉ1B��h���#�^��o��TX!�L�j�W�1	��
��:��e���"�0�H'(����Y\KP��+�(��w�)(=-ٟ�P¥U�m���b����]�ټp������|�j����Ҍ̵�ag�z�%6��G�&-o5��Ԓu[ܾǎf�����W7,�ӕ��f�R�_����
y�'U�/��ˍ��j����oJf}A����$��&@R'���T�n���+34[EIK���J��-E��\*��o+�������배'#�������9��K_�W,ki���3�۸r�ƾo��{Nܕ�-��0آ�(K}�
R�5L���eKe�W�L=��4L_��O����fCe�������3M�6��Ws+)�_�Xyϴ�%nh�-u������D��?2�	����Q&��y�{�rs��t����&{�|�o�(�ݱ�8�m�?<9��xq�sV(h}҆?�;�2ͽ$L�33�9@��:�|�`����rĝ�S�	�ǜ�hAV���">y�@\���!�%��W?�+���	�I��N�K��r4�����#ӌkA�6p
$��R��=�`��a�$Q�����"�"���u��`���z8M	��u��W(�����{E�n�Z���N�J�ˎj�����`	9a�(ժN)�����*<4!�S���D��&���ٽ�̭�`�b)�{S{Y��N�X"!}$�-��wV}YǰD�{S�ͅQ4q�W�8*�&O$Qێ��½U7�+�dp�Y�-( ���������,��\��m)���j����w~]z;��e���w/� �,�(��md}��N�&��o��sg�� ח�2�~Y�y
s��gX��je�ϴ/��k��v.�TT�j�@�>r�B�?7�t��������:��V�I��]�1ޫE�b �͍����cMw1��m�Q��-�h�〉�,~ADɂ�ߺ��+11��Z �y*�� Of�e1����Է���N��������:� ��� ��p�����#�Co�.ԫ�=�T�6�i��	(��[k�Z&�����
�|s�, W�iU��r�Y��}�&㌹�[n��`%MI�`=�����m3�U\�lJ���|~��b��A�)�#� �n�P)���;t�F�I@7j���%�x�AZq�k�p4�%��ƿA~�֟��T7��ꏅf�w� ����/DcTlj@��f�-����
~���+۠
�{gxF8����gb�h���g�C5N��R!�
����C�C��� ��݀������?�=�2ni(8IѦ�\�[��� F�
I*����������C�?|���@Y�U�8��uHk3�_��N�Y���e�e��E�0J���{�[3�U1 ��2���Z�
��xw��_d�t�b�@7�j���7�`ʣ
ʗ`���6�XGIF�����@ɎU0aoϞ^��u�h�S�x�� �a�b`H=3�k�sG��	L���;���l�5u���غv)���� ���Ji�����W�p�&D�>l<H�V`t���d�d{�ǅ�I/�)�(t����Q�¤���ΰ�u_8��NbU��ȣ�k:[�y�Wm`@�X �����d ����쏍{43L�E�u�<����Nr"�t=���"Ey�Z3P-��=q��_�*����������M��"�U�P��O�w�f������/u�RFт-x�ڤny)�Ufb�?�c��<��f�N��w����E�ƺ�������g�v5���Q�5�Ƙ�� ��@m^,#W�8�c��&B��|��%�n8���t����O�
�]g*�Z֬��Z	��C ��*��yξ�s�`���+��C,��0'����.g� �_�f7\�'�S���t��f>7W�2���2 aS1}}+H�^x�'�]z�_t�t��Yjͩ�ۿ�v��_?#-(���3gz���E&�k������QU0n��~nK4����^����uK7Y�T���ղ�/9v3j� ɹN ��S
n��g	F]��Oc�B �Dke���X�,�W���d9�36w��e%i�M�5�C��4�Q���ųJD�()j�Quٸrsj��̛}��������Ćо�g<�e��1�)V��C��ke�R���a*�a�}o"�^F}����4Y�Je8���@?-��7|�^������F��oH������ӿvEN��'t?���jrJ ���LT���jeF�Y��Y0��?cPr�W��\v������l	�}x����J�\�������^�~o9�|��}* ��������y�^;yah����Z�_h:S�R13����ݣ{��S���>��-�	3��G��j�L����̫�s1=���}�K Ϙ=T���t䯒�"n��B�
-��e��~��s��6}*�
���d�)˽�a'm�$>�+^GD��C�N�Ձ�/�c��2�	8�B8����-霉XPA�y�-�P�=i2��]�Աǭ~���K\kt�G3^�O�
��e�|�R9�q�T���ݽɒ��r���J�Q�V�Κ&u�jrH�]��jt��O��֮���L�T>�M��4�Fv��$K%M}����!>��ƛ*�0w슬��a�)J=و����@�q�ɥ�@<�^Wz�Ϧ4�5NW�<71Ơ�RmI<��[�k���b(���@q�}|��8�&C�c^�>3R�빞jd��mN�}����# ��۾_ѭ�؜��Ƚp�$�Q�?>od��ʚMz�C����$2�`�rA_���Z����p������~my��m�쟿��'XT��^c�3%�?z�,�:�CY9@?M�CS�[7T#�@iZ��c��C��vS���v nr*m:�J
 ��=�s J�����*?��ϜME��~+4^'h��/��8��>�|@/���qS��:2��E<bg����"���Z�5���b\i���37}aw@`��R��"�,�R��y)�	��4�#���1�[jE�J1ڛ�{�-�𴯯�O�Akm����ڄ�w�/�K�g!��2ߜJ5�}����-�Z��C�ѿ�[>Pa��y��K��.��ps�«}���5����u?1�1��S��l��&w���~����{��4j:�f�I�x��ev<���;�.T*	���_
���Lߊ )�tʲ���yM(D�t�$M�<e�H��ؤ�ͷ�_�y����;D��_ �����t�_��\��}�w5(T�SO��bH�Mk�� '��8'�M�J ���U�����J5�yw7�H�!�a�Q��,�̤O�p�]�E�^��\ޯ���d�a()�^"!�^v��� ϻEn�^Ϯ�����y�4LT��9՘�;�6��/2o���һF�f`E]���K6���A2��@&r3����JaF-@�%���������H� ��z{�s�v+��%	R 1��{����g\�CSSo�C�h%!Bz�f ����E����(\߄I�<��3��P+n+����T!g��WB��2- �ͯ�>��]G�ƭ�ը�P?�`)�ǣ؋tE�["ń
`x)�_��$��ME��>S>�:�ð��Nwۂ;����{淗�#6������G��L@i����7�{�T�m��d�}�C��8YMw.���d�T���� U��
��������:�7�-l�_�ս�&S�j|��B�w�
.�*�ꨴ_��m0FE`��W��o��W3�RWj��ރ�T����'L%��ΰ"��ali�I�o��8%�h4 �L��sI��(��d�'�K�]�x��`Cm��!���V�N��4moY��d4Y��^��-�A?Há���9����>+|6m�.����H�Q+�Jm���,X����X��w�/�eZz�����)������R�ث��dS*��^�	���8F��q�R!�O����\7�}쑟�}Y6 �6�}u768'�K�bނ'Q�j4�ڙ*��Jt����g�e&�>A(��aW�޻8��"?�h��9�B́�{IZ����K(��O�o�苑��u������ͷՑ�G&BM��=�lզ�1���0_񱣸��W��W�a �Y�gh�d��i��1Qo#
�۠��������HÚ���Cx�����n�HQ^���hM5@����X��FN�W5d��tnG ς���#��$�O��7%���'����)s�b���!��f\��0]�A�-˛?ZI��bݮ�K���C���7�(a��?�|#��jO�ǫ}�p����� QD�?��o}��S�ܾʥ��UVG�y�*OL�o�X����]�IQ����H!1�T֛�iL*S6@�xbQ
TZm����V�61鿹�b\y"��&��0T⋽� G�U��^����呂�E��� SA4��ĉxxڬ�7=	�I�����j?T�藬!�`���:g�S��-��)�9L~��� H ��$t�H� ��@�H�������z�t�qF����/�my/-���*�:���S�}�=N��'*x�����ь�K6^:�}��o)<a�_8�'�z���hX'�O�q?�r���#�&=�����o�;�/�W�RU�䡛���롍
A;�L{?�\�2K���PRR�w����s�� {��!���R���7��A�S�է����hUsi��w�&__U;��C�6��%-��O}vu�9q��S�f����������� ^�5⏬���&�z��%�8��l�3�K�5~��`�	�f6�H�fW�ȟ~M�H*��mcMu?Q�V�!Y��d��5�I�tp~%��,����Y�gB�0_>��t�]����ւ:O���J���T�uTT��=>��(��4���H���Cw��)(�)����%�Cא�H������k���5.�̽�<�~���9g<�S�|P	i����!�tHw�$�M�y���1��f���[��$JN�ޙ�)H�~%8c9<�s����0Y�j=���%���ɷ��"��U�(�Y:
z5}���Kj�����jZJ� SXz%�U-VhI����3+�5.D��G�I�D��Y:Rl?)m��k���;��	w�Hk��>�����u�aD�,y��,�� `x^�^&����7C�!]��+G�bH�m�`E_;��j��ύ|}fa���wD��O!'c����Qw<3с����h����R��﫣2xE����AhJ�e���_�в��J~z�"�'o���͗�~�@�>b^jg���84�����s(Ƙ�	��T��M����#���X$.�3[��������ܖ�S�'4�މ�6l)�HQr�
�����1Be��]�ݔ�[>�ۑ�Q��Dh����6��<���RU�oy���a��85��H*}�+�@y�&�*g:#]'�n<��iw��~]<�g<>��"e����Z~���o����x��Q��TFN��-�����.�ȭ����L�ˉ ���tI|���]�!!��C{[|���&F��W�	���.�m����[fo�^���<؈\�g���|�ga@��g*�r�'/����]�sF:1;CN������
���JO*Oܠ5nd��6��劁���ɜ3�4�.���`�3��w�L�����܁�	��3�(�kG˻�ytb��s`i���V1:�v0�[�P�7��U��c�T���d�?�����^@��X���4gs�����3��RR��\�����o�+�ʢBWOy������5%RDF���Q�Y�A�V�<(�N���#����Q�0�չ	� Nr'�Z��3Yb��OM����%L♓�Usk�����f(忛��TS��M��[=�w�?3�������_�x�l}��ݒ�����H�M��_�_n^O�OI��M��D=�k�fR���K�]�h���fݦ�`�s�8�C���~��4jD,� h��7$�\��u�dg���a������t%.J�/w���9�(#W�\�F��bm�MPJ�`ة�c��'�'3�e����Kw_v�M?,��3C-���1y]�xY����~�n�J�|FL��=
vݮ�&e�/��)�C�V�g�
{"H�a��w��2͂>�MV��::�%�����&8����·�Q�z������ܐ������wl�����|��cZ��rvhk���L;�S�q�(�T̐�ꭝ��'i�\m@$s�	�7�tϟ��qd=�3�~Е������6{uٽu%א���ZA$Y�\{u6R��S�^���~�i6M�#f�y�!e���wYaL%{z�c͵`��.rj9��ir�S9J7�<p/��^��0�F��i��H�3��g�tO8����G�	q�eC������S�����r�B�,O���2BOп@E���J�^�0�j�w(�X�R�V7m=D~���S���L�i�����h�شD���j��h��1�u���P� /q-����v{��)��h��rG����Mb�E�i���8W�o�Ј���O?u'���=^���/��!�%�a�������rx$	�=����r\f~O�Q�~ck���:��\
/�}��n�-�ɼG,�R�w�Ǣ�p�\TP���c�3���Tݐ��������=y����|^�`�x�ZkĒ�;��>j�k\�;>2� N=�y���苧�!d(OK�+�����;�M�"ڸ���C����1�_���DМK�<	%����s
��a��2��߳v�{�y���xؾ��d�~0cROZ�ӴN�i
+X����Cx<�D..�J��(��7� �:���J�+��c4�+�����J봓g��v#e��t�U맏<�ᷲ���6����-�5;6W�Q���)4dgp���5�΁�Et�Y�܄�����*�hа#g���tnQj[O���]��fvY����H��#mm3<U�K<�s�ng1���cn�wk,9��C�X?���~��K�a/�W���EO]�EzojɟG��~_��h�"��@WC���,�������%Z,�9)ɂVFy���Y�[!�=�(�}?���z��tjQ��J����~��5�5�~�EN񥮰�A��Ŏb�/l^�MΗ�w�lxOJ~Gm� b�)�q�_�=�4K��1*�!e�B�K�'��i`�.�q`��y[��Q8C��،�'�V�}
*�|Պ�[}�������S��К&#I��%����*�K�6��o�E+fn8���s|�F��r@,�d�}���_p��F�fH�,��q����k9�C�HwX�O��4�tC����7���W.�q~
9�e��gzi������	kT�7!�U�N>�ǟ-��AfzQ/u�^��6_`�_���dZ�� ��_CrCADwy��<��<kcdl��V��U��/~Z���o���$*r֋�������Z�Bd�o�o�-l��	���w/���s{f:Ѿ��´>��B�����2��K~���@ �ȵP"J��Ժ�-ϩR��!kv݆�H�l�T���n$ö��)������&T!���X�V���k�#:![�qO� 1�@.���c��T��KJ.���1�l�`�wW���k_�bاݰ�zW5$ˢj\�qm�m�����<�ܔ�w���WR� 	���iN��7l�2�k3�Y�S"�[���_�@���k�B3�S{K�r�`k�@�0M�/jkS>�Ǖ���azY1l�7Y俩˫]��m���1=}��� ��m�P�+*
옰d���I�޴���m��u�`R�K��.u2p��jW@Q~��wz�]�u3�e��jc@\Y��6��<+]q�<N�U�Y�H�m�~��J�����5�E�����8�-f(�;�%�I��(R=6�4[>��q*�'#�o/�﫡�J��g7��(^�΁�l�+kX�N�^��T�K��ի��u�R�IA�qE.P:i���3QG�q8���)�6�M��<�E+�Z�5$�X]�--7�Zر�������[3tB��ǋ^��#b K�{c�e�{�u0)�'��v������-����5�������6e�����K֎��켹ї{0?)]Hk�����uZ?����Ɯ[?�sh��z7��Y�vYܐ�N�.�ʂ5���}�n���2 -9�t��zր̅J���9!tdE`}�]e	E�˃��"�VL7��Zm�HzZN�f�WWH=�����~������l��Z�`�����#En뮤���/_K��t�0X��ƕ��`�pM�!�J�:ԩOf�F֠�8&�nD�V��#K޹�Ρ7�����m"�Zb5��EhnC�J	[O�e�:E�M{�2�?#����}c��:�	z+� G�����U�?���@I�s6���>;3�W=�u���$d8����L�c\�i��[���M��hw��ܣ�s����'�>Hp�����y�O
��+[���d���q�7�A���:fP�/�{􀮯�|,��%k��f8��d����.��8!���ۘA���,D��q��f(�� z4Gր-T���V�� DY�lB}9�por��Qt!@^�g�b6��f ~��&֜��P�5E�_�Vh(@��/���X��W�iv�n/�a�q���%9H�����,���~������˳�ź�YJ�8M0�g��ǀ��iE�&�f����f�OJ���A�����ĵ�>�z�J�c�Y3��*S@l{�>�g��K�s-�)���T_[WI���k�b��w5��:�vG+P57�:�6�ŔZ����Nkⴼ2"$�ER,7v�+�5�"�I��8����N���!u��yEk��WO������?��}oO�|;�<)�w����9��� �������n%.���)aI��~�D�$�#�Ks�����$��ë~F���5���#>�>n�h�)9@ҙ�ȓ[�feH*�ZN0� >��
A�4œ2^���o��N.��Gj�a�b]�@�5��iύk[�̆��r���ٯI��i�CT�hw<�T{B�P�Qq�����FHԺ�Ȃے3�wR\ .�ص��a�J���Xi��緥`��;���8��j�ђ��I?l	�]��w~�����<�ne�&�� �!�g�!r��
���U[�r�[.�5�X�\� ��:QD�C}-oNd.���A��9��%|8q�h���H���c���8e�B�Gd��<w��4ˀ+���ۊX�>鱥�~�W���QZ��b�
��4�O�ͯ+WI���a�.�ٍW.R�悻l딫#Cy�]�{ö1"d�xD ��c�LMAn��R���#
?��*8L��QC=��峇*&�pq*�y��U���&f�Ja2�{9g�}:w�Ѥ2���}���k�� >�c��2�?/��;�P�[��|^L	�hX�~��n�
�����'���t���i���ؠ��%o�s∽G�m6�*Y >�_ym��a7+�E��!	]��婾m�:�.K����
_S߲��'}}\��NR?�{�.v@M]����U��_n��D?b{�����YZm�U��2|�A�`Y�к&�dӞ��S�%W�oW!��ׁ�Hl�\��Ť e��CuV��R����s��q�]��A�8f��M�$��[��J���ot֌�+-oʹ�X��.}�^�x}ڍ��ߙQ���sM(�9W����y���S��:�w�N�DG��x��]ih@O?h�����#���5��G J�t�i{���~�v$i�\x���}�~C��
`K�16��g/�#�;!����ߓ����~������K�f��{B|�qh�k�/��
�3οκ ��2r� ]�+�0D�������S83����C�~n�?p�)��M<ǟ��u�A�¦��ـ	9���fm�f��+��`�%��Ȏ�o�}����D�^�#b?|�J~�DK�������ʆ�s��*�8���p�;�Y���zKg� ��w�������!`��!���t����0��b�oi���	Yڜ^��&�*�Π ��]z�؇u*�bf�����-�!��Ƚz�RP_�#�vG��Hw�������ŗKd�֬#j���'l�d�z�hH�g���|%�.&î�������zU�/d�t��F6=�+2�v	�⽪�JQ���[�vP��q�_����_�[~"��>oSRf�T��]��\��p�$'_	�HYJ�W\Qq��^����m�r:횚j�À���&vJ~<\~���pm�J`y�RSvODV�-���:oI���(�a�7�Zk�"7X�}�~��Ś�~�8��m���/��y��E]ӗc��C6�����M0��ع�Q��{��V1E_2�\�x�&�L�޻����grzz�Hâ�^�c��L��MN�%�p�@4^�*������D�{AT]%l�M#I�U�/^/O�óY�� i0�s��9�b�: H����2<�����F�j���H����і�"��͛�y��_��\� ���ϡ��\��e���5qh8�B���Y�	/�RxA�E]�/պ���W�E�L\D�V�T<6��GH�>��öXd����S͍�~��|��W����yK�^(T���L٥}];��g�6x�g��W���p���x�|��#�C@6�J�g�uS8z�=��m��}����,�G���$�<����{��J����$�_��)]/m��p	�.��z^�٦Z�PK������,��h�U�T~ɐg>!3����`��o��U&aK�v�\Z�,l岼5�^���*O�Aqq)i�߆l)�nV�"��x�kK*�YX�tã��F���������l�.����d��������^��~|����4��@��)2Q�����T3K��H�<�z�h����ߒ����KTr[qﾝ�]w���!?�-& /���ۿx^xn��S�a���p "՛��H�p�P�XDvZ[��d��[��*�]*������^�����7��8��#�B6}x��e_u��l�>K��?��-��g3�%P�o�]�7o�n�qgt��Ҡr*�[	UH"#K9�wLWx�ȼS����RΏ}��\w��:QͯE�����K{���$M��ȣ�Ջ������gU�(r�Z��lf���j=ʚ�2�s��#��ق�F�W�~.v�ڑ8�?L?����.8�:0D#�.��Q��$NY��O8���"7�'d�*��HVY?Uʒ�4k)7�9�Q���p�}�2�M/ ٷ��N��R�}l���!X����}�gp���aỸ�_���)WW��z/��ڀ"NH�<�C�7lFn5|�\ɍmmGq��8��N��%��i�U}V�L���|���sW��6�����݃t�~o�P�o����/�`~�-c��:I��$8��y"B��5��M�8����	�y9Ҷ�l[��ÃR|���z��4�񹽐��1oaB_إ�P��\�I�\O!�2"�w���Nr��-��,۟_�6ŻX��C��.��/����B��KK/��}v.�3��8���H��FҠ󍰾?f���}m�ێp�4��/�:P��w�F.�!;����P@��";���r1����˝�blt���f��a�3��3!ELŌ�(� @�~�&��렿q���&�q�9�i�ܴ��V�-���LnO^[�"b#���a�ڣ�	�� ��^{�A�_�PJ����g��R��B��M�֞Y[� �W��q6��+
�+�0�����P����������M ���֯W6��p����<*�^�dT	�A�H�F��PY����G��^�=⣜{�d���AV�Q�c~��u����b`��C��B��J4�"#�C�h��$���_��uV%���^�!v�'�?ЈpD�]Sԓ��jj��Y�!+�[���c�����طSY��0���6��5
��v[)���x���?�;MM��w���V����$I�Wd�O�?��8�!�����uk
N ��H���G�Y��-�xdwP$-��2�|l�����o�¥?�x
��\�HAEֹ&�vw��:_+�Dd����e��v~��P�o"�����é&_�B���~��N'LO*�֠$����8����_�]*�4�������YE�%O�f���7�jB�n2)^�Ԣ�!�?��z��Mt���j�cO#���D�Ǆ��}�}�����3�9��()�|i�}|������݆�N�fL����X/7�������??m9t����Mm��1~���9�򸲜Ԃ/f��-�jTz7J��{,X�[|�xQx�&��߽̓u[�{�_�S��z��}�p�����p6IW\��#6���߻��p�������г�F��wx*�/W������nY�����ag��/��z�WH����Bz���r�t��KY���pM�|���r�!��v�\��;���`�qn�K�yP�>�{:����3=�"L����M*����_c.�u����WK>z���K����zӗ<J�Ǒ.!m�S�����f���]���K��%�4ץ���w�U��ly�)��k��C��n��8��c)s{�=C���!G罭/BQ���w�����d��k�w,+d��N��h{u��v���	�V��Eӎ��f2�?���R&��3�B=���BV��ǧ0������Cu���v�3�ip5z�n�Q�$���C]0��X���̍����nđ��9�'�Ւ�e���7I�H�`,�=`�Z��?}N��V��3�9��um�
�"K�*Me!�q�잆�m'͇"���s�Ƹ�:\2]���x^�0��aw7A���:ڟӟ�rYq��K��CU���L��5\)�s��\h^���I��J����Q\a^����`��y3�+8NL`3k��hX=Y"�T>\|�	]�mG�:�ͩlE��4�1/AF���0v�ѝZ#ڠ�z*k��[�`Ζ���RZ�{�:Z9��;�%��!����L�RU�D���g󝉫g�S����P��զ[��Ǧ��6`�6�;�֔�԰��-V��g�4(
�*�5�c�T:z�y&�����O��ҭY6#k�GzZU�{��� �@g�cs܎�KJs�P�����U0n~�^$��#Y��:E��;�����*g�x�%G�S񐉆��)�5Ƈک��%�[f��o�e��-��VW�[x
�3�'_vY��T<���,�F��2_�R'o��$Sl`����s��r�`/�O��7:8),°���#��׆�{�"^~P����*j�Q�ꩦ�I�+!���P�wW���t%��Ab�j�!����#R7�͆T�z>>P�����I����\^V
�Z���;�R[�!֩W�w񇳝�����+��g2�b�};�7�"�&��
%��u^Ql/�����LՅ��~��1Trs�����E|OK]�	�1z8gZ�ʔj���K�E#���wc�/�k
S�Z*�|_�{�����Z�{Θ7 "�/��e�9吕���ul^\HK�C��&h+�W�+�o�Jr��\O3jĸI��{h�Y���'��l��P4\K���\�>G�a�[5���=��/����-΅�9k�io�E#��j7��w�_O���̽%���u�!��( Ѝ��p�[�׆~�@z��;�6EC�2r�?>UԜ� RV�6�?����Y�tO�E�-X����̱s��ϪX�b�@
�J��f��P�G���99&�l +�IYd�+�zZ�_�y���/�$o�t~kB>�R?��d&SKQQ��X��E�U�� ��ѥ1��5xٹ�p:�s��|���Bx�)y�L�����sQ�sp)ǻwb�R�3da���R�0�i�:O�s��4�Z)�Dr�����D�B[�/l
���杧�����P@>�J_�3�M�JJ� %60�/a���|���s�n) n:�+~�u�G ����O���k�⴯�p�((�l����6��?F�����B��g*�=�Akdr�^ ���^��|Xp�V�K~;.ּ�P"9`�s@==��~�D���u2�Ձ�3��P-����c�+����{yY������f�c9[�C,m['�ˌoۗ5z�/�����p0�<D=�j�*�է�μG�!ok��t��Y�l:jd�M��E��P=��`^r�E��8�C��0��z��Aϓ��5/ޟ���'�������| ��Y���#�Y���W#l'+Q����zy����n��i��.���8��Tr�Q�E�^+�
�@/���nWrug�T�W�Jl��c�Z��a���b8ln%�p��^DO��y�t͓�Om����\��Z'6ئ��o�<����8���\���x+Lݷ"���0����8��7����:�]�"�C��s�t���j'�1��R�5ڌ��EV,�4������0�]���]3q*S³�w���~��n�����Ğq��C�ݻ��>{���}��Bfs��}��Dd8�:�B�r�ڒ	���	F��]y�p	��z�i��8�����;x!�I��0�i�R�iQq����M���1���h���qI�A�4(�)�$���2& A��q;�|��9�a��9N��\�53W�/W��u��O��/~q$E�d�/M4;.����?�ˈ�� �=���ѿ��P��%�&�����f�4�18���)8���𓛸��MhI���q�w�Zlf��:^G�j�k�[�R�������+��ݝޓ%5�A��S	���y;n�;Y�r�E�9�!'�g}Ь,
q#���Z��w�����Ku�(겎$��٘��i{Dj�s&�'�k���?�w��:drA*5,� �nj:6_����@�B��N�y���S\��jT�������b.��2��c�q׶qv]!h����"uѤ]۹���Z5Zy���z%��_�����y�����9�6����#�1d<m��f*��� 'u{ �Xim��:�WC�h���d���P%Z��W��Ω�+}���YdE�E��l����V*�ߵ!�O����ӥ�K>���I���M#��hrs}�{��y.����W�M��O3=U$Dy}r٤�b���K��r�ёf2���c�G�\jэv�b�Β��"Ɉy(���+_R�]��1�H"�J�ڙ"v�|!�Dv�Q)e�?��y���IS'J�ܣc�j	�4N�Ms��;z�-q�8mA�࢖�͊��iÇ�L��7�W�ٞp�r̕�{ԛdP���Sa�̕'�pb��������]��s��=-P7���x	3�RLޓ�~���8���V��7L$�{�5Ar5A2���m�m�Faɀ0�*��ń2��	�K�'��3W���|�iqQ �&AgAA������d��.��X�R��4Z>&�|H�E�]�4ᙫ�tV@��^8.�NWq;�"^�����u�TI�k9`�n��!�g.�w�����I+X:V!0�-,H��Qq���S���+s�V�Ã�P��Z����wS�[�HX^a�
�_��ʝW���UY(��{6Y�����Ib|wf?����t���ތ��&���V��~	�����1�q�C|�0�"jC��UZ� 	K�)��ջ8���_����5�W���\��xi��ӺMB�G���v���	Έ��p��B,ȕ��@���N6f������}�h�k����Ǩ�ȢDΰ�b�`��[g������l��e�R�M��#���x������X���U��v{(�ڤ��=+W�u&\�w���QBh��d���CY�Fo�ͦ]<��=��N���,�q�;STa���y�s������J�I�4Y2OG%����/l,^�Z�^���2¿�1���«��h��6����>��l�l�gk^?�Xi��]�4�Jߛ��5�9?o� ���H���װ|�����jN꛵s�S$'!�[C�0D?��M�&3�J�(��8>��u���z.9���4G�d<�%CN���sXA�QPTV�g!
Gn���1�ż��r�C�����=�\��:瓺:iP���O������g���_��3�ӿ�zv�s}�VR�v�"�Q;Onj�T�Q1X ���� !�sxA�Md:nF����Ռ�R�Z)��}ﶴ���
��\��a�,EO>ਇ�*W&�{sz�B?���R��6c3���I�z�bu7Y�������t���Uq�Q��Ϫ�������YK����"�|2VA��� ڊ�6l���+�-v��o���0���A��}�A���ڕ�o\#=R���7��I�R� o�.h��2�<����$=�u�\���6����?��yoT���h\&_v�E�a3}�X���}55���T��u�Itˬ6I��}�h�~�3�%S����f�;j�����ٕ�qi��;��fm��_e��^��7�&��[�w�Hί5���}�����̕z�,Y��ci����8�Xÿ��莖p4�L{Vn�v������s�%pnB!:T(����f�np�FR��<�G���kX6�((g�'�����:���� ��ԁ WS�[[���h��a�;P�����_�вZ�B"oB��F�5��c���װ�c�݇l͈�X7>����8�ȁ�R�q�C������f�[��k���ˆ�8Q�z��rh;�eB��	�a:ڳ�F;7�.���>g����ןo�^C�l���v�`ZT�,	^��qǌ[bV��C�;١9�qlU����k\�$�ԇe����Ҕ��ԧW�
յ<���ff��<t��7�����C5����PS��wz�!*ULOg��,`p��޻��n����3�t��q~�y����׈����lYR�]\u���k� �VL��j� N��` �a���f.1�[�{C}#�����v���ʧ�a�@���k"Uo��A�8���ݜ��)��a���x%�	�IJ+�Y��Cx��z8�	�Qa�N ��¥�Vj�[O�e�-��8�6I�f	ѥ��g~��W�	X1���|$3�w�U�Ң1�#6�1j�1�q$=WRd$��0!9����V|��6? +�M�3�~z���ܥ6�>�5V����vW՛��C�)"�%bv��LPQ��[��J֤m�m�J���Ŋ��&�B}��UUV,E���]�s���0罾�����6Fb����+|Py}AT4p�9���'�����jP����+R�ˢ�?w������FK��lA&�dB���ɕ� �U���`����A��Ӈ�	�[K�����';f�-���Ũ���zf�h�Z�ߒ=�a4���uu�螯���D�cM�{��X����,��K���	�DƞPY_<q�ZP��]H�hߍ���%r44^�-����r�����Wvl�1Q2�5�O���K�X��}�|��E�
�]9�*~�;�/m$A�ܯ�s��|ٴ��Z�iP�Ϙ:�_�n�^e���j�����ݾ	�n�9]�MZs�y/�P��B[��l�0��`G���ӊS�W�-˒�
ş�Y@.6I'��A�FO�څ��^���T� �`�}I.]z�/(�����^Y���p�y"��u��P��~+�c%è
y�`� }�5tBs�L�#]@IӰ�����Q�&,�#�_2:nL����<ޅ�U�N��Y�~��!ω��@���c��4��.e~����`�]������������*���X4��K��on8�7<���6��'X����ԯ��߱�b?�6H�=�+�e#��btZN2��:�o[�����c�e4���f��9������zK�s�D/N�&dń�Kl=N
D�θ�7y]����.K�1k��r��b��^��i93��Xu��c��%b�0��M���ulr���!��|� QPXV|�j"Ӎ��`��^�4�)Y��L��O������\K��g�a,N �_�=�Ҷ����:�='v��VՃ���`�e|����&$d�质g�F�kf�<���8b^h����I.wJoѸ�D`~��[���������R�=N��uehi���9CR�0��I�2�w�^�X3�Y�m�	�/�\f�(����,�)/u��=���E�!�]�|��ޤ�_�Z�]�V3Z����Ia�a����^��g*�g\m'תP)yqO.���Z[k=�����S��ʅ���J���}��.��]�'�����z�ᬜ����G%���D���o����Sd3����2�"�9J�/e|��s���B2�z9���.p��X�E��ak� ϯ,Ȣ�������,����Bo�R��o8>��6�^��^��\�A�
3�}}�rYru)��<�Ru���s�i#A�~S�W�I��!b��������Z��+���� P����;w9��b�>F�Ŝ&i^�����W��e^���4�?�m-�-��[�r0k�ab�ޢ
�������G�'X��d�� et~��H��+2���i��D�ؐ��>3g�H>�G �۝ȓH����򍚻�D��ovR{���dֲ�bbB+���ԑ��24�À���7�,?W�7�+�,@�O���2v؟���ǎ�i��.������j7:|zH��H?�ܻc�=�2^�7X�K�;�qL��ʭ�z�G�ʧ��[��Wg1J��  ��-0��uI_������h�b�4�m� �ђ�cu�qi��ca��������j�S�O_p71�r/�1�x��m�"��7=G��,؎UK���]>C�y�~Ó���_N�w���2Om1@ A�v��gn�怄�>�h0��4ZB�%eK� i`'|Z�E��qL�[� � ���^9>�m�[�G���y�`��k��Ak��)���*YO_ �fw��)/{�y	�H��Mt<s��&�?�4~��.p��挅nL��̾�����1]R+ ��^ �n@y����Y���'v�=_��@kx�|R�Au���L�nqt����p��E����ppS �?|��,��}���
��XM���QT����_qB��1��:��5u>�ۀ��?�B�t�#;��
tM95@��'U�V�i:=�ٲ����6K�t�E��Fh�N��6K��ȳz�6���x7k'q�������D�K/��h �F�%�#_K�M�3R�0m��$�0�'���ɂ��2�E����@!F�8W���<u�w��lK#��	��[큇@��� vW 벒:��n����c�)A��g�O3��[���́�@68y�=�53�(��( R��B��m��dq]�on����z�p����C)9�Y��l��Z{`�f�{�[X�Fj��@��;D\�*vЁ�RH�����O؎� ��΋������}`V�FR	J�P@ ��Q���Y+z����c�h�# ΍�q	��i�\D�	zz��	�`�bH
�y��~إm��!�FA�#�\X�~�D!��,�T�tf�{C�@���������Q 2�p����q]5"һ1]jl���W%�x#��G�bRvì�U|�q<ewv;3�O�=�� ����.�VL�a��M�b��jl�X��Ѐ�l��9�`>�r�R�Ka�fh���1r*T=s^��"���I� �:퇨���T/Yp�s$3���\H]��N��J��s����v����J��>�>F�c��2�z��?�ktúK>6��tO��Gpw����c�zΐ�>6�|���@�奚�Ά�������+�w�D5?�s�\�� �p,]�IF	�Ë9��UxR-����{ CJ���,�[FO�Ѐ�}���I �4\��l��8�w�"�$nX���;�	4d,�V�z7^��M+M#d�zn��I�Pr��t}����BP� ��(˜�F� �x��d�+����t������כ"��<�f"�5]/'s �5E�D�������ɑ0��=�5?Y^����" (��|��|�LC�0 ���r�G_z�*��"��"���Td���F���].-����~w�W�! ���C�jFZ<�FJ������M�ο�&���P��N@zJ�^�Nz��Ao���6!ۼ^����!)��m�fd{����4��?�j��}�HWEG�?
�I�5��ij �~� >u���Ew��^6��uq�B���`�e��"��7s���>�x� .�ר�� )R����B��$��>"Ý� 0��Cl�E�_�������j��9�C%E��Ay0ɛ>ϫa�f�4R�*m5n�E)�o8�dV�1��i�ŷL~u>�0AQo�Sp�5�����&����?Uz]�������z:�E���os�)�q�/ ����b���s0S���ķ!o�ؒ���`:ɇ�ڲ�@x�E�~vW��Ğ5���u�-Iy����xa��Z	u�Q�����2;U�ƕ�����g���U��YK�k����+��RϬ��'�?[�l��"�>��N<�'��J}3�8��"#��N��!k�+��_���Ɓ�5=;�7q.��Gu�Y�N?�<� >�S����/4�;�cu4�\yY�C�� sK��+i\�BF���W͡���%�=�#��K�4ӡ
����`*���$�3 �_2��Je���C
M�s蛐l�g�ygV
�����O6$�ӑ���&�3DWxN��:a*���!�`>�b�!��A�@���&���饏�?w��0t&o���"� �3�|��%�~G9D�P�d��;�9�� ���k��U���	�`������ޛMG��y��F ��j�t!e�t||ɳ��@a U�Ò��!��/�l} IWے�3*w�Cj��ϫ���'�9Z���� ]}�nMm�/Q��9�5:�n&�LESAr�4�����mFރ&�N�V���P���|��=���}�']��W$
���]��%��"��cb��J�Wc���)�����GVKv�I:��Q�<�C�O�������p�l����0+�3�[��9�35�M�!W��M���-v$�d,���@?�"���$/��A�I�� ���@���0��Ϲ������y�A�N�������J��$`nѪvs��g��=)E����|R�B�񚷄ֵ��:�'�Y�C噸�-d7�|�� ����.��5�(/�+��I��}�?���|'p1�Z�l�n��q�<�����������z����6ʹ)%�.���j�+��5�&6q*�C����=[��))vP۝�Ԕ٢�n�}$<�ʘخ�"���~��ν��۽Iw� 	P�K��{]x�H��*��2$	���#	���l95/�L���Q���݂�`��^��D���@ <��[�v�qWGj��*IK���@����\���� ���h���nYЎxx���(L�xĳX�k"�
�ÏHYb�~�d|��ë�F�5�	�!��Bˠ�S`}+ W�������$��R�b� Ȁ!G�N�k5R�wZWZ�g_X����ٺ��_L��V�;!�/A�f&��_.���xjٛH̀<��ǃІ�b�^���8��S�q�����O�
�!7q^��S��~}|���ϒ����v�_^^��w��@N����'������>��+?�I��j7��/NV@꫻fѕ7ϒ��R/o�z�{ZV� �h} ���\���Yc8�d\{jTN+Kmӻ$���"�=uc|�\ 5�ӻ-�xg����ߞ@�m�*=���$�\vv%5�� I�O��	g ���y�8��"�??m�d��7R�� �wmj�C�ȿ*Ŗ�Q=yc;��@�a�KwqL���
�e=�Ժ��C��j�;z[�X�$�%!B}�S��-  �.0z�a�.f =��^��-�4�B���Y��_�j����v&Xaxg�{�k��mz�.����߼�Sz��4�5^�e�N��|
����[��%/���������*{�w���k�
�J�()��+!5H7(�t��*J0��%H��H݃�������/�%��<����9�:v�
�E>��`��:�|p��񫺋�'��k|jK�=A�tx0�Y���~b��^*jZ�CSS�G�6�/֊ 5A"�CM��Mc&U�<tϗk4�Rs��z|�d�^,�G�?
��zَ��G,�q��8�6칥)�6V.�[%�F�\����[�@X��*�իk(��k��R�}p� 9aTH��о��R�x���b���ܱ
�0�ڗ�Ap�q�7/�fN=ɍ2��3�<�
:Cb_(�]H@�{%�J8k���$� ��B��+�����\��ҵ����|Ќ̚����a	���/g��٬/L����K���M^�Ҵ�E㬢����!hy��V��������rїpr,7O���rj*�� ���7�Mg��8�4fK�4�׌�/����]Ys��$[[ȹ��+w����\.	*g����Y�ad��	k���B������A��~����.�F�K�U"���6J�ɥ�h���,��+[ˏ� w�D���k�y����0���Y��9�� 4o�
�Hb�z�<�PZe[S��F�4�%��k3�i=���l�`#�h 2ܵ&U�3=�����Yz��4�Ȏ���X��E"%TDn�yN�l��-���d�"G{0��W��'������4��@8�ö�"/��i�FJ�h�x���=rTp�h�Z�Z)�)i������}0� RW4�L��?J)���4��U�����(�B�)Z�Z�`$^7�i�	R������4w�~�"s:\���-���[��g��Y���K�{J�����1���7��]�ӊ;ߓ\s�tp$!o�ǵ΍1n�*�mEB��#�^�ڐ2*�q9�[PA��a�U-�-Jq�k}��,�cڻI�p��a��A�ݥ�7�k�2.��܀��z���t�e�x�h�u���J�,(X@�?#:�o=�\{�*�.��ʲ�D����T�`����̷����)���w?��kqK<u�dF�0M�<O��pd��S��چ^���A?����s���է]m��{��&,j���>�Hnj�(J>\-�|g�tt	�w��:���U�0������"���B_���n{��<5����'�ٵ$��yy��F�+��}u�����6��3���@��`rz,_��yf��P=0`X]��kj��Z��V���O�k�#P�j�e+9�.b�Ƞ����L���Z���9��|�tS���(��4cLO��9��?�*�mE-�ѹ���B�j|���`��a�1y��ޱ9���^�sVj;ƺ��|P�Z�,/�т['�?�P�V)�L�U��I�Z7�jsX	k� ^�{]\���	/���p�#X��>[�������6]"��`�������g�T����{���G���kn���3�ס3[�����继>���ꖥ3�1&zYS�J���&�OL�s�-*��0�S��Tp����`��#���o�j�Y:��x-2�����w��#"�����nj��b�uf�������9�J�w�.��x�Wzf����&��Zu���竤w.�a^�i����ବ�N�xs.��9��E��k�Zڙ4�l ���>�"
�xz
>@�Z��Øp�,���l◡����^ʠ�,\�e�uǶ�Mw� im�$��?@�_@,�w7RF|(��	��I�����|O�0:y8ͱ2��ri=2lg�6��s�����!�k;� gQ��T|�v��We��h�[�j�C��k����*�����D�D��ރ�*�q��
�UN�nh����
JP��̾{}�����"�j��s����-�vZ,-���Qj��_g�=ƞ���(�=��{#:��*�O�4��I�:P&v͡���\�	!~�7M�%V�R�V�!����_lL�nӲ[���S�~2ʲ���+�����#l?V��Y��{\4s�Zr���$S2��H����ܹ���r��>�����ˏ5��F��r�����i:*��bCu�-�L$��:��,���{�}Ò�����H�������Xz0�C1*�3��|(~w�����T��d;�'$|��6|�w��6�#Ԋ|hC��AW<k�hxt�exjnlڴ=M�]7j�
K���.?�ئ�:������v����pc.sG,��ˎ���>��Y��)q�`#S{�ڳ"V����/y0�j��f�?aZ�Щ�S�c 9��X����gǦUhGd�yi6�
��]��{_��f�zT�����0��m�{y�o	ݧ�%ʡe�zD�j��r���m�l�����|}�_x�gN&�C������RV��J������I����R�<j�{�J�R�s����U��Z~�QJ�����+槗!�����V-b�JqRt�C���Y��I������8���<q���B�䨶>.�|oR��Y��8��Ak��H�m&�qK=fم�3��B[}��*2n!`n�����ݳ)�H�C���`�57٥][dK��I��p�]�3��}A��_Ѝ����CA���'�o�}8��{���SM��֡�	�3��y��܇�WI�]����
u�'�V
���U��@��9�z>�g�|�#C��b���Cg�2V~�
�W����s>�h��-�Hya�����j,����1�˅#o��6{\j�Oi}k�d���7{��wk���Q���-���W���.~�e���G��<H(����c� Q�����6׳�7�5g�Mrᗐ���)�ΚZa��VVr@�?h���]�V^eG����-s�8�m׀p��ܻwf�K���&��H���Q8h�2=���R��g�˰�n�%�)ei�0�	�Mk�g����^>m{ѧJi}�l~f��9�} t�o�<�7d(�A?�t%>��T'z��kk4�g�P4V.5L��jt��{�Y}Re����%p�D���v��a���S7F71ez�E��?�5��ԩ���,�@�����s��^��+�o�\E�38�H\����*4��T����]\4Z���(�W�݀��e@����zf�s��ɦ��r��s^ �=n��<H��T��>�C�]��ċf�����L����f�Lx�=@��F�䠌�j�ϣ��q}��f�_$�]c�.�]H ���}�G� �\���n����R���Ʒ�	��]}�[��w{��Q9�ܴ��u�ɼ�d�jAq�%I��H�)���L�Ύ�e=��c-����v�ԺTB�s7F���[Gߺ�G"��jUX�??*��f������G�i�8Ӄ�߄j��^��T{�pԝVUN��JP����C�R-�����6�@�h@�Uv���C�@Xٹ�1��4)g�q��q�Ƈ��4D1��)��}S|;L��S�9�%��Fd2P��d�lX�N�2J����W�CUuD�L�B{��0릳��*kN)�J����T�Na=/���q��g9O��D���؞�[^$�^����?طW�m> �O�#ӥ*`�4�8@ٌx��x�Rlz�T���W��w������9�,����M �x���<���I�ra+y]��8�,�hf��<�Io��K�0{#��H"��J��)��8m~qe�l(�gt�C@i e=X$�ּ��~-��%6��'��IQ�l���&�h�&6����@�a�Zɨ��)�h{�Q���k!/5�U�h�*>'i/��i���PΞ6��<��X�o��f	�j��x��`v��Qϝp�I�l�re�aݸ��,l�-��]�����YI�Myǟ��l߷7�!����ߠ�3��R�Te/��D=Fw���G���׊��?�71�U���dܿޞ�Yɇ���߃j�g2P����M���y\1���՜�&K�ϝ/�1�I���A�Y��� �?k���7?������sv�XkFL[j�8���H͗�r�L�{߹�܎Ԫ/��ą����C^-#��g��eC�暄#�xD��ӭ��63��5�Sj�����#/�~�ٯ�����D�yAm�8�WCV0�[P�)��2��= �њ�(��U��(�U�jX�t����"♍_�9q���1��_ź��/�|��җ�A��!�[D��\�W=&`<�Jƹ������U"0�����s�9�^�t��O�j��A�-W�@�WA�C�F9;��h
�9��Aw�5nb��q����-kL|s�F1���N��u��_ډ8=���*���N\nL�pZm�^����b%���wz��������l�,�e��{>2 2�q"|h�O��t.�8��>2����}��g�.��;�-�cX}�3��<�`ڞ����^��V-�M=���������u�lsai@�݆T�p�]�?�L�,f;}��q�G�H@�cx��'��1�M�=�il3�i ���4�>ȬG���37w鐜.̓Q΂��})6w^�B)<|��Ш�k�co�mD�<��:�����ix���-$�u��w-�m�|�6J�*�i+�����`;�G%����BH�â�IӋ�Ui5���[*�%���?pf���w�K�m�o�aijB��9�N!z�V��D���U�<���]����#?���>;2�����'�>̹��j�}bͼÇQ�g�y�I�ӬrIx�򠥛\@s��5��P����~���!w��1<�Q��ۧ�s��E��<�!էz������L�v�/�J�h��bHz��W^�ėO~"��-�x����}�z��)@hҎG�WU�WӬ5���T�
�t��a��LE�9\�z�K @+�!Wi����X&�uB�.�,�����^$-SpW�0���/��rN��G2�ʤX��M=`����I_K���P�,����ї�"��q�x;k%[������	/�{��}Br{d���a(�W{_R�oI�%p��Q�ha}����W<cF-��o�֖O\+���X�� ��L���;QD�?���r�R��~����n4J$>')m��ָ�
��"���R��z���t��|��"vYH�Y�q@��`͕9���a����}����L�B��02�t坧���E���%�;J��(�|n	�j���L��Ŀ�Q]<}�Q�_�g�9��"�L��ۗ�E�v�,�F#�e��a���.����]��̩�03]8|�є%;̈́��,Dl����)&{[=hҖ���|����3��nSƈ��ѐviqm~���6*Dw�#ˑ�uN���݊�Ѧ�>Xً�5�c�`n2N�����~��h�iO@�mo�~w�odӯ���w>IQ�faJL���N�MRw��8+Pwڽ#��������G� )�H�Lpɮ�p�].ݝ,A����]����E�+;ϋ\:k�z����7=��,�X��#���J�^�%Y���R���Ƈ�#�����w�f�I����%
	�+6{û�/h���.��f]w�r����۵��A��O�6y�,�V��}૭Uu��n��˃o���5Ɖre��>���@tJ/z&tkÛ<Q���ׂ6�r�g6L�[�p�t[��Q�![Kns�kSsy����Px�W��p{�E}���_�7�B�͛3�㚑G��zE, E�(�Ŗ할]qX8�&�Ś�C��oc�}������ƁC�̟3;��W��	W�����0XB^�+��Ha-�h�m����9��c��{�uǆm�Q��<P��mV9����a�U�d\Ha��K�'y͎����k���p�#�dѮ'�h�xS�����n�h7}�¾�_�����rX\���8縔\�{����iףyö˂��Wo�������BSE�\����y�d��Z�wt��:��HX�T������U�\k��j?��$J�t��������a��++@攒���CZ1��wd����ut�o��I�<���@f5�#��#{?D��RÞ�#�C��%'�-�l^7��M匡�����s_���y�$s�Ný�ll�!�vrsC�I�������ҦέE�.9ϩ!b��
R�Ҡ��G#��A����Y�|��s����UlT$�R�~�
Gx�
?���]^�}0�;�X�����&Clo��^s�Vd�91'[׽���B�7o����W�{[y(�nT_��Ơ[���p�a|3^AxlXׅٴ�}>�y1����z]N��j�@�4�3��ǂ�<�J�� ���:�5�Ҧ����Ш�[�&"J�z����!�	M?�=xKJo�C>��Q2�u̾�b�6�_�X���3��J^xoȎ�t�pużC�H�&m8�
mM��[;i}m���
k8R��'���zo"��Xv�h���VN����:9�K��%�|���ڛ��(�)��r6�`��W�-�8E+�_!6��gX0=�5EV�1�Ey�v��G:~��Kǵ*�TԞ��哸bDz��tBn��~�vwկ��1�Z�<�ʲB~�n��`|��Y$���%���=����}sF�NgA�?h��V�
�V߇�,L��f�|���t��̕����4!�s!��ȅ�<�d�Eڴ���PFO�׌�'Ǻ�i�YT�s#ji}lȯCV�+�n[|��'���
#+^,U�!8���
7T��3���./�?��\#�t��j�������;��,)���r�M��m̱��q�q��)�6I�#I[6�I:�=נq��۽+*$Յ��N�_�:G"�Zz�/��b��h����D�X�1Wۂ�1�<>�ї��7Y�=O�}���Ǌ��Ő��+�ߓ9�
O a��m�0Ye��Mwu�j\���t�%��,���?_�c�T�۵���m�1��������$��K�%�����g>r��ba�(q��,�U����u��w�?�le��I^�z%��y����q7��h�2��t�}9~S�}�!CT�ɳ-���M�j�^׎6|lg�wpj�4�(�R6�2)�֦q>>w�X}��OҰ��Z�S)��zT$l;�^��j��^*U��Jf3�,P��Ũ����euv�Ѹ�&�
�4�?�Q��Q�ub���G�g��q
�HN�������}���QoNg�����\�h��:.����#�$dbatn��3�j*D�(�O��uW0L�X�if<����8�g�n!��e, Y��o�b�j]����O�􈣮}=B��(8tj��j�b����$�Q�0�Y����\Ͽ<n�ɱW����P�W��O|�P���ycd7�݅sl,gk<E���4<���/IE��\bL��(�
h	$��+�v'�'�Cs�="������R2-5�G�n�M��Թda�͡�6R���ֺj	�6��z���C���%3i�n���&s���gN-�.���|MG�y������,�q[3�5t�q�G���4�LY�`H,�,�GV�u�Ů)�;?8b�^zMG��'�#�l���e1T�v�$�#K���������4�4����ʕ���Ԣ'�b�<=gr���>��l]�ܪW�ͥg�n��,.D��1$ ͪ��_��� 7��;��u��.U}mb!���#���'?�@cJ�u]�������A�<G��5H��N��Pv8�ܶ���c��'��֦D�?{nu�P ���^@��&�>�F���4�B\̊��.��.P��c��� �{����H]޲�E^�r_�(_ɝ7 ��5e�H������<�A���B`"�|���'J��K��yDӶ����Ӿ3�r{�r:��zP���w
Bq�v@L�����\����+b؎��?J���[�1붐�cv���[���[����Pq�Q#����fO`���I��ԡ�y)��Z�+n�C�������v�?�L�ӣ��cs��=���e9�$�o��3u���e�[�k�mb;�D�?��2�o��gcc91nv�Co$��/�L;��l
�z2uW~��߼Ƚ�nj���0�#���kM�@p�����덋�!D 0���@U$5iM���p�9����F&�(��|}���m����k�6-�|g��0nٓ��opl�ҏ y~H���)���X\����%z(݋��)D�z�����և����nw�b���⻿�!k	i�.��:��m��o x�I��-'���.�݅��M���mE19��IkL���=I������}���5?��zl݇������;[���?u CX�����FrN+}�K]�i��27�$X���@ ��u��:/w��C�)�)�M@�R7|o9 f?ݏ��;���p�`S��=�.x,ys�RQ´�c��sF�i�u�d��hm<&Y������Ë���y����޲C�����c�f+P6�*�nP������8���\�[�Ƕ����P��b�"n�T�̐&�h=��L�gk�%�녛�%������}�M(��}�H��A�IҴP�9ⴆ2t:�I\�hgXE�a�1�\��,��.�����@��qW+_)o	O������<"��C�G���=�|�W��� 1�I�A���W���<�Կ��G���3�k�q+�C�"$�\��}���q6��ƫ�2eZ������$U��������N�h��V��b���E��Q������;��œFW�8��7�"VkĂB����"u*��2C$`�f㉜������б�V�����>�gD��M��)�+��_�3}����,�PS�Q�t%W�
�J�����S�4�5�%4!2[4�/�H�7�����ך�bb��q�B,ح����W�41��: �@a�w�RW��M��Y���U`�K������O�sW5@�<g�ܴ߹��[��pm a'�O�ʗ�������[�����{}b��߄B��%�x�# ��[��ܢ�Q��|����A�M��C�KI�I���Eoi��Wc���@�	�	���A�Dw��F���(�)'kw��zD-�2B��r1�f�Ŗ[˔���ku�I�P\{��/�^㩮yׇ����m=�X�7�x|}��^v:��Y�=`�SeHP��~z~���2ғ�d�'6��b43���ڜVZzm�ߎA��lH���S���;�q�$A��LF���J�=���t���O�����! ��Ѱ���h��L ��[�s)�����viM p����ޖe�PKc{��T�p�%y��@hl��(�ʻ�%Ξ�uܩ�Bb��*�daR{ ����Y����ԽS�)'����a7=���qCu{�}�=L���f�g�	�����11��	�e�j�fGc�KöhA�*\~�k�#C��b�K_#�s|Yf��I�E���c.g��3���GօS���{HEi�16�UP�L��XV?Y��X���4����d67���hC�H��%!4����m�!D^�D�h��tA@/>� MW$�7'V���\w�?�N���}�70���բ��+�<��0yl^����W�I�*ګqu�b�^,%4�ᦕ��FKG��V��֭�d�we�>J*���5��Rɥ� �K����V�T�.�9Mf��hv4@m���w�ED���O*�l^7V����{(|�Bj�ܺzms��sT
�)��E�l�L�Q�A�b��F�[�l�,���EPx�>1��,�u	5$9��!�.+Qϲ6�Q���qΘ�L���-���*AU2y*�B흳<���] �C��~��1PANf�����O�ev�ϭe�����u�>�O�H�׿o����Z�� ��.$���s���a�P8����"A~� g��P��<�_�s"9u�Fupp[l�	io�z�d��'^�I�t[?�iw֯�*���AA�4��(G<5%�Uj�*|�P�������M_��wB�����^�?QbPy+I9g0=�\�����,b��E^'JP����ڽ��rĮ�n��]8��j�t�g�U���˂���{_���a T�%��Z��3��������ҕ��� ̻����٫B/���\���0��P�q���3��� ���Խ/6�UÎ�%�2` g盘�����L�D�z��Ǎ�D|k�m�Osc"z~D��,���M��5AU6^X0������@�r��!Ǉ=*d>�$��_}1��z!���b�[�e)2ۃ�h�F$D���th��ك~����������RE��
�,����ER�"�=�=׶��Z�((7�����ܰ^>̓�l��nAn�h�n'NJa�Z�M 9��(5�F}�Ġ�����I�Vbe5�J�v7'{�a|Y}+�S_�)�D��j2�p�F�åK�������������4 �4d�9������h�/!�!m�lp,R��{jR&�H�!3!w�f�:X�9�;R��~���>��:O#�|9�
�����z|�\,��8Q�L���m���3���tIQO�D���p^a��}<R�z�É�C|��
���w��G�t
��|�[���tN�6> �����j��&7��6��!��+����s?E���p��W:97�]��E�z
K���yc�X�C�l�e<j8~����b\�E���<eK�Q,�ȢO	����}��kٛ~+�ز{�O�삲M���� |@=]a[���C�vleޗ%�~�*"ZK�*����R7  8�kR�|�Y��ʯ���Dc��ʰ��|F6�$[>]����l�:D�,�u� �4���ll�	�I!z�M�@�d��`(aY�=1��A�PT8�*(k�^�V�W �
H�T���8뭝�M_��Mz��|C�[�ʶ�֒Ĩ��g!;�7�;�WY>Uc**��+o�
�w�[�n�lΝ�|�]�Ѽ���34A0���5�����}��3�ZQ�OY5��ˮ�����9��f�
�V
V?Y|ZB��LE�pCR�4y\�E�3�/�N~&�%2.���UW͢Nf��"(~ ;�0��-x�q��
Қ1R�z�ix�pܡ������c�%�C��!Pf�Ӣ��v�̭[� ��������zD�;潄C�MP��uleB�7�E��/u�u�I vh�<v�hL�������
������\���և��b1bE�ۭ�F��<E���o�14y������Y4j]���QTN+N�Ya�߰�6A@�odRְ�I�� Pa:��)�x��6����&D�} ��	E����}�:}��gn��M�tQ�J]�T���������qq�i�� �e���Y�4]�U��,T��R�R�F"�Ʉ�ܐ�_�8��y��GyF�	� ���* X�ᴣ.�c[{o�g���E��]��܌տ7/�9��X�V�l�,ѭZ�ף���EKyP�ۺ��2�����-�[T�f�M�O�:�V}�{���i��������7�-���r<��|�&W^@��d��BC��U���!�֚��ؘ��I�n�S���ɺC_��8��QlT�,TT�ڃ��zG���\ֲ)J��1����J�v���'i!�9�l�c>or�X൛�6����MU^��A���dW�QE���3e�3S�n ��	N6�� n�(ġ�G��{��_J��8+�<D
AY��/�
�na\�Z�e{���?N'�#��<~��//p��Vp/�y��:5������ὴ�8��EM%z���j��\� w��t�6��J�PD�Ҽ�B鯱gYφ ��M{���q��Z.���b�V��(��ڷ��Ӭ�6��hh���=U"�f*,���6����O�I~����?��<���_�	�h�[d�wb;�D��J	������u5��P��M��w�~m~A^C�NQe��,s��^T�?�Ǣ����o�x�1c
�����Zw�a�hk�q����Q�=Ӿ�U�v�LB���������i��<N�2�ô�-m��_m=�!�l���x2�Iqbv��20}�b6s�yƺ�y�w�u{�;���<q��eP�a�~I۪?w^=W�������Y�Q�H�In@r��-��|&���~2�l��4'ws�}�t�p;�'V�0)H`�@Fޘ�6�{u��-X,����6��$��
����>��鷋0h�G��T��_��°݆�E�n\a� ����Mt����Gڥ�;@M
{�f�f!�M�q��}w�f<��@0�u��7�����Ow�A�p�l���tDC; �i���Wڃ�%{29 ��{�� p��)9%��N����c,�
��B
L_]�0�6Ӆ����y�,"��OR�)]dn�ǬY�����5�i!?Dʾ��+: ��Y�� ���!�.��珢��6�����"ڗ;שs4��	��}YO_����4��!�"p/]��AW̺!Q8�����DWD�$3�}� ���%���t���E'��#}`��\���;��-��l.ˮU%���R���	B6���c��;�ڊ{H��IXЬ(�Ӽ���.3VM�v�&��I*��4��OO���+�9u��F�2�J/��!/�����n� I(�f@��i�'�j�Hw���y�A���C7V��*���YU�>����=��=>��AM�� p���e�ݮ�͒��ڔ>��;�BFBH,Җ�>E������%�����}+���M%�*X{^��OJ��`(�tu=��e���tW6���}$J�(�܁� dm5����	Z��	�����e[Մ?O�r���
��(�X��\��zH��?D=����O��zg��� <��Fj	�O�|�"G½HK�>�`�9�Ib���^9�]�^�ih�/d�F�q�ۏ�n�JL��uK�1���ʦ��b���Ni������EƫOZ<�����F"ό��p�]b���%����K���K���]�{�ƣ�U\�u=��1���K*��N]J)3	e]���ruƌs���s߸F��[���R2e[��äV�۔���;D۪�6@�)g�X��8�w�R2R�g��4t&N^UyJ�{ZBQW�*���K��5�}s�+�AS+��a	R5J��%e���D�݂ΈR����F���i��&l�d��z+Ñ�&�M89�9�e4�{(#�.	A�w���R�
TM-TU��T�6��_��k�K}9�/:f1�l�J�
�K�a�_�a3P��`g�A����W�s)��4`E�K�ܒ��ӭ����ɝ��97�
?I"�ԙ�(��R�v�����a)<�\��m㭗-ꋘR�έf���Z�wN-jo��PiD����f?�tGd+,�]Fm�"�C�W�ȹq��?�#��r��yu
���M��%���-y���gN����2��;7�u+;ݏ���C�)����W��,��.G���Y��a)��Mg-�ǌ9s�e�ˮ�x��p���3�����4+ݮ�F�>�N���wN�VFrY�Ԗ �MO�G>�lWm���� �� �f��?Y\�$��#�;��^��Jբ��	�O&�V
�7�R�O�	����E|̯i�z#hN莨ߍ�l]��ޜ���'��5�-����C@¶#%� �:�AVF��b�&+���w�y����҉�52�0:R���/�dX$�P4X�P�`x�6�z���ɮ!�U��L��_m=��I��!�Lym?\�ǂt��#]3�J���	��*y�3K�~���r@.>�'�>��k���k[��O�gȗp�O�)r�d������K/�j*�Y��|�����N����|^ʑ�#�.(�.G��Sc�L��r�`��3ZE�{�3T��_~'C�#�'���A��g559���-����Cֶ�7;��h� �v�� c��b���a�:ؒn	{�m��?�=<<��v=�V��d"ԩ�$������p�0��ɣdr1r���?d����		#D�G����wr��a�f�3ϝ�y�I6J���o�����U�'�I&�?4.>�&�4����7r��{nÊ�}��,�a�Z�� R�Kڨ0�����n��{u�#�j�D:8���Q-Y�z/���sz5%��i�+Y�Dh��oKJ����Sz�D�1{��/x��r��b�%�C�V��-�p?�,�F��!�߶II�e�=�߹���
xg��/-��Иl���N�����ɡd���s��kUx��PS2��7��h��?<�t�)}f�!��8�6g�5*���i'�n\}|Nvr2!��?s��h�C��������xv�z�WP�`}⪩���[>��b[�Q��+>WU���2��t��{&/T^�KsR�$P�n���X�>2d�_j��Xʴ�����̡ȳw�ېV��T���	��۞ԉF��ɅO_��X�?�$��mTR��Θ|����Uv"i|�pb:/����t�C�ϕΜ�T���	Ee��	���r��-� �/��E ���M�D�GϱwOՅ�N�l^�#`EZy�I��:)y�R�o'uy�;�N_��b$��r6dS����ۢ<6�O�X��2�7R���ρ��������J�ss����!qH��6>U�ɷ��%F6�-vR��X�*�t�*�0��Q0%�D=������.P�����^�w�*��2�
*�e9�1���2��%2�)sW*}�����Ry�5�T���7����m�%Ӷ9�v�����̉7Be����N3�S��F<M���F�%Y	1�Ł�LYO���;ysȢuק���Y�R�CyN[���oFy(ֻ�Ԕ�<���
,��[���滐3XF3�5nfe��F]qZ>/ {V�?��T��,yy'p�Y�����L��d_�D����K�?��l�3T�xDj�锕�L-��E�?��<�V>ן��m�ԭ�k�qZ�D����
's������;�[m2�;s�a[b/||��
D�4�^�����yˤ���_�yW�"k���PB{����ͺ�hXϴ���*�FU"|��oR~����~68ՂZ����i)t�7��f���~�T��<�����}�	�X�i��ÏvE����7K���idmo���⬪fKd]ѭ����Tmm���|�E��?�����ҏ���'�Y"��Z�w�\�1�����Y�]�d�e�xB�;�^խ9
��D����7!�O�d9���4�j��u��9���oŖgk�fXh�KrV(R�߾�F%"��JԸ���0����N�TF�����,�;.%�=`�����3y��j�X9ʮT.E2�%%�����q)�@�K���|].��^�
z=̋�KA���J�/�S���C
�@��m^�hm �h~+�_�s�!�ؖ��P�MQW�oY�Y�/J|��\�/4�hx&,�E;�����*҃[)��c�\��0�����z��\S�������?KE�ī�	ʮ��ؙ���K�.o:�}2� 
��#�}�2OutN�BW�%�������;[�Z�U�o��k���j�"�� o������<�X�r�����wF�Z4V���[��á�q�ؕ�-4�tJ�;+�؄(���$B�~��Nm�Gct������መ��h�r~pLM�`M%6.K:��X���F#Yn�lXkx�D�����nn�r`�+C��9{�.@C7��*���LKQ-�yԙIc��(�y�w�y�~���1��Ē#��b`�c�tc���>���Ѣ�A5��g���JH������ٟ�>��jM��(N�$���lu����	�K��u:�-{X-OjE��pbၩ�ce_N[������9�"vk�,y�i"AQ6r�����2-W�j��F�J�l��W	��?DN�Z�?5Y
R��/���ʪ����u�"���
RuJ¼�"ʔ�
��H��:�-wZ����1�<�Q���M!�b�"w铸~�Z�.��ߞ��/���ѷ����*���gk?��61���.>�~��K>�^�|���WB"'��RWi5��i	&i��)yDCHEWH�K9��7��ȫ�<��V�h�q��]M�G(�!�����7Ϩ�3��Fz��
�(	.|�~���c��Y�m��{ܷ`F�?��z�B� �z	Mb31x��s5��*Oc�|�sK��@��WR~Ց���|ߙ��I;*�ܮ�$��/�>�s'��*����-�^���G��m�J�-�}�����t�*�n�����v��i����ɥ���V�_o�J���pR�\v0CMQ�x��%&9&n��:���c�X}4�*��!������_Ӿ�Y䜡��jR�62O7õ� `�M���Ε�e+��vj���2�����^�{�b�uR��e�n-$�&��-�
�?t$XVf�C�k�K�+�G;�fpm<�e��Q��{9͈�"k􂬸j���ްu�1�F\]p_N��rF��q*�.�r�Y��.�s��`e\kՋH�{7P[.�V��ԁE������C�k[tYa=b�s���T��ﲵ�:�|���}+���/�e�'숷V-K�5o�`ظ�W��XK��F͙<9��H�{�?Ru�@2�x,��{�T����Y�b�!�J�ǃ���uֻ;���OKWv�ss�sd��-_�����$!��m��S�;��������Dpmg�\ĵu�]�{�ח����Ù�*�V�s߿{ԕ�:J[a�Q����!_��V�+�οE�8����E@q��n�g����\U�����&�Oо.;}��Ʊ�m}���o���gv�O;�y��9fW���W�X/�bu!={�{���H#-�3�e׹��ø�+B���U��~K�\E��u�s:�Y�'e��s�I�a=2d�"����0K�i� ��q�.˪ i��-R�O{�'o�y��^x˜٭y�O�_g]I_��z�b�+:Z�;hy�'m"�g��FD��+ьؽ��I��O��Mw/�J��
|-����5l���yI�����tӖ-����Z��T���aI�f`��g_tt�N2�̾�ZSƎ�?�	Yt��z/�Qe>��b��٦w8���C͙�[�-��n�Oz�	���X�C$SD��A;��_��.�̬lX���L��)<$���f�,���t�/�;j_�}7f��߲}���9����W�`��|ΡEu�S/� �`��c�U��A�bQ>��6�-���-B�z�o�Pʇ����+g�w8�o�7��<G����?�a�E�ĵ����Yҗ�%�+'QM;��ʣ]׸���ԣ�2���(/FX]�R*�zf�,���G�Z��sn���'B����V�>�搴O�/+3����%I'�w/�ED�L}�.�y�Q��=��||�8���jFcqE�܃MS�>IJk�����̫����
��FL�"��vS�V̺�r�-
���3�KD��Y�.m>c�`ZCM���X�� ωΫ�yb!bC}��!�յ��8�켏�H(��4���Y�=���pV_�zee�7�l*x
WB���@(���?����s���o���B��5/e��:rժ�˖�n`��e����&���^C˼��5��rϕĹؤ�Ï��?�j���[v���w�_�6���F&�্�E��rT����h�zZ�0a��=���n�i�ڪ���Kx���O��l��皅�%��3�5����������`��s��A[��X�	c�e1�9.��
�/��E��J�����`�v%!�}�L�Q�]�B��r�6������Uw������Q��hΛ<LB�{��GG+
��(Úә<Cm��j��=�7Fe�������j��Ml����s���H�,�,ɚt^����aQ�]ۃ���-*H+
H+ݠt�]*�94 �5Hw%C*��94�ߞ�}��x�����^׊s��\�x|�b-԰�7P�SK��ju3V�_�D��v�ǭoB�{��ů��c����Y�.Z�7�!���F�j����d��r��~����Hq�򑸸���&�f��u]����m#jN�Is5��S��R�7��L>�O�����w�Y_�2nF�q��/|#��]�K�!�+H����ڎO�-�����H"���ϗ^������Lx_�|ҥ�2��������`�l��
����Ս$>`������|��q�Bcu԰���]/�{�،�BG��$�Ƅ*�8���eH!�ז��q1�+��8F��z������'�w�F*��"I�9D���M'i��)e̤��Hܣ*J �֥�}�o����������l�����N\�1�ARnPM�}p��Ҁ���I��|�B`,#�8��<!j	`�g��
e1df ���J�N\����Ё�o����ZP��=,�Z�B,6� ��,��G��>2��&�F�t�Z�֚5�ҥ��M�ZUl4v�������j��k�$�8�H!�a�iޭGg�R�x������+�}��fedj�mF��u��|�rq�7�J�9܄c8)���u0�.i�"�<}fM#��C|� -��e#r�)��[������Su�g��n�o��N�d��R�R�jX�Xgg�0҅w�g�^{�����wi�5�{Z�־��EѪ}��0g0�l([��|g�EG���u���l\)�ʑ�:��r��'�qQ�	nM����{���IsW���B{+��ܞ�J�K�Ano����2�Fʐ9���f�! .�3w������,)�1v56U^گ	^'���Wx��c�w���=��U�dy�k�]R�y!C(>�C?71���c4vP�t��{�����c��m�������	a��&�O+h��T^.2_{�;��j���&|	���C���m������֬�U������s�=>i}�^��J�������)(X�P��r)�@}]����X�y':7�lP�ܬ4���"3h/ꖂw�Jx_/R�x��2R4�%���
BC��p�D_CP�aG[�!t'ld��,vס�4��z�߄E�'��Tc��1�CW#B��@j���N���zM��M��ff6={3�O���V�ޮ1�;@��]�QU�q_�#i�M,(����?��o>K���B��ۨ�&�"q��e�x��:�H6��z2&��&����(@㦚���i�z��A�Q��b?�8����_Rɡ�"��Ź��wXك���#T�2IEU"��s?���V����@B�9X��Iˬz�%T�� �c��i�Q��Re�x�˃�v];�@t�i*��\�tU6ͮ���5�����Q����������� qe�{�'��vh�?�W*[i�z�v�~$��j�� �_#�#=�33:ȵ�W�'�i��:�j����@]sL��Mm���4�:�ڢ�(J�$n±|>/�,�"��J�!�}(lt�w�1ԛ�F���7��=�n�xY��K�5�c(��YŒ��ٛR�� ��G��P�r!����O�v}���2a���y0����� *����Y�ڐ�i��$����Ħ�p���U�Y <v�x`�D�Y@�nJ�Չ"��8l��G�	�$�]]SVR��DmP#�q� #�˖_��r�@�+uM���2�Q�44��LH���G�6��Q0Ϩ�L�B.ĝ��ߍ�b��X���s!��`���Kp�e)�Cz�l�̸�˫^��dVz�r���!$�#$�����k5���E�`���>��1���|��G���i�П��I��j�%k�ʁh�x *�:�����Bü�U��������l{�h��xf�hޒPtfY�3vEh�="Wo���a�:׆����Zl9����8�>�J�Z��m�[�r�����TY@���Db6ʳ*��(�R��	\�u�4�K�ƳHV2�t� �E8�Z�uT��B˟�~ҟ��7HC��7���~A��.�2�$��F��Ifw`��k���h��+��1���ˮ�cD�ܝ��)�Dt0y~�v/�k=�,.y���}�B�����\�k�I:s���X4S�����z�/��	�-�?�.�?����%�6��
T2�%�'�4���J����o����`3=�y�yC'K�o'�����߮��P��/#�Ɩ�,R�M6W��)���'\��rԠ?=��%r�ɱ~�_?��v���qބ;6�&��w׀�G�t;��~�Ѭ7 u.���EHv��i�S˫����=^!�[�v$6����^�_:N �1�����]O���Ҙ��I�)g���/�HxI���ѩlg&��ǐ������~r�/ɂ���Ҷ��\Dd��c���<~L��
�0G8+N"K��W��$"~f����Ђ�/7"��D��l]�I�a�L��s�f��Ǝ�����xJ��!I�N�=�}aCA��q�ǥi[�R&�U�0!�"���~� p�ب<���
����ir�	�p!G�N1����6��{��!����R�&����ˉ��۰��G��F���15�##��|�з��m�� P\��R-�`ܞ���?�Y�1���eV��T��
׽�ODp7i$��q��AΦL�tM��Cz���H܍�n�"��c�鹦{vcD�̥�0a]+� �M 7�3sXX>����s
�����qoX����,��S�]B@���p8-�9���:���xo�s�F�{bK�g6@�p'��Ў�.>��?��$8�ё��F���B$N�P�·���o�v�f���]����:�U��ݞ���C�K��ε�!V������Q��<�w�G��q���{J� ��i�%�M��Z�j>�4X:ow�b��/X�CP�?ӟ���o����M1�������������{����;�#W�*w�3��x>��3��� x�&����a����/��Z��9׌�%�=�1"��H��|�u�S`�ߠ�!>�X�wQzSw9Dۧ��{��5$q6y:���\wA����we� �.��٥��/�~+�FP����-�j�Nfr����:��Lp�q�1*�ώ	�o��Q��&1m�i��~��eW?�����0#��jA��%�oU�N�� ��}��k�9k��g�ט?����Y@��k(.+v���I�i�Ƕ���DA2@�� ���4��E.
H����G|s@�{��9�eG�\����	�3kT�L}��XW4�na9����;���8��:a����զOVN
0x0S���@�xU�oTFX�6�Ȅs�Uq����'=)�Ɔ����=c8��pH�u�� W.���^�\��Ƨ�ILW����\�H���es��Wpx_�@4�R���
dJb�\�������IVp�p?�ְ&@��Y6Kj(���6g��	�b۟�>���X��L� �nf)���v���6��[����lY�x�k�3G.ɦ\�=�࣭�Ll?�� K�͢
��I�m}���?r�NT
�S0s�̳}�����8*��HRQ�نl�]k�mJ�Q� ���w<��7��������ɋ*�<y���[&k�gE�g�ɇ[{�	u;
�D5�]��:'�� �t�Q5�ʇ�O��P�+��Wr��;�]�T*cD�li��X�)�۟'�����a�.Qnt��Â{ѕc�7q��KO����`�;�]��Ӟ�����28ٟB������w��15�+�)b���@qLZ��ION����)���Y̈��l�~�m�
6��+��s�f(<Ȑ_`F�:PbG�q�;ޭ��Ii�(���x0 F
��� S���]A	��	R/ `��{������]'0���02ՆIzV��vS�\����	{.j�*����dP�P���JK%\h�������r��M�3�oH����J;�$�C5 �o?:��2��<�e֙������sk^gk���w挞?�n����������e�bb��1
��^ m�?�"���ۙE��D- ��l�{Y�2phx���eL!c<P&�>�����G�� #����F0��}&[!���hl5 �v�F�,:z��]��}�kNem���}�MM�9���L�؛�cJE����������v���������gM7��Y�%����W�k�,E�H�e5j�x���
6?��ߥ^Ti�������V�F�հz�|���I=�Z�4b�&� k��&<r]ߥ�����й��	@F��+Ϧ}�Հ$�C#�F���l΍��Cr�pS[78j���5a��οh����� T�.䯶SS�ƨ�/f'1jb+����0���Sz�հ�?�Z@����{��J�Ȓ+�H\��O��엢X�V���KPK�#���rޑ� �qW�����6���F�����\�Y]����,G��C-���#"5@����Z`�*D y�r|v��^�S�o�	�ΫO��N��B% ;<�@�p���j,��Y!���{�����1�1�/����V�*��m�Ll^l����_�n��m&��5'X��>c�ܤ�G�h�W����"�XW�Z#Z� ��?Ru#~?��9���!"�y�ra2���i;|�;ke���S�	$:c���]��̡��|���whAB��{��ƆLH^��K:0k���P�����m����3}8��%y3� �[|��_�3|!��]�hi4V��Lɟ���a�v��$n�]Ǧ�+d�\�Y��W�y\�����|Q-~/F�%��n�������ˀP_�Ϲ-��M���-]^��Y�'v���~>f�r�j�BpG!5��.�-JX�t�����S�>�$U��s]z��{�V��gd�
,EJu���m�	I�w��xD0�MB�������M������&\g�\�]��r�I�O��~=���/����A��.E���L+�Wa��E��(n��m�4���|��gυ�e�)�M������"&����z4 �d���$�?��sn���<��uX�T�q)'�o�<!�Ax|��^T�h��l9�j�������y��M�~����mn=�����ϲRf0s`���NW���ށ���|�`�R ��xz�\�8���	z�c��kI@;r��<��[���ܕ_-�
�M����A���[��**`�=��YA�W�@2�aي��,p���Xp�
§��k�x� ��=�YE���o�Ub���,�}�*W�*�)>#r�rP|.���\����`�V���e���o����ԑ��f���V.:��B��mǡ�q[E� ��E���\�������{\�q�~Rȳxr�f-���|̍v4͑?��	)@.[*�e'�%�8*��Yrs�K��)�͐��3x9���*�HF����:�Jc�"ru��r6�V���{�'s~��+��43�&0���l�㔠{і&����wҢ���˶��l�;p�l�~n(���JZ��%.��-�*b��d�Z�ڣ�!��J@UJV�]7v���+{��xEY�4�*�K�}9u��B�Z�^y�̋ �'��a�$����a��}EN��粦{6C8k�����	�v�m镔����O�,D_T躘ϊ�\�)Ff�k�6�v���H��g��� :�M����D��]s�MN�!>:�*5���`Z�xW��;�У��u���I��Utѣazn/���u(>q�kl��:;M"��q�=	X���{i��qw'կ�����-:�q�痁�E'k�M��QGEq�t�<_�`J3��5	j_�>-�]t%��F`Z�~̱4Kh� ��V�Ǿ��e�ƾ3�ݱ�¸�y=������t��5���:�|��s�5Ҏ��ڢ�5���.)Ώ�nӭS����j��A::܇�|��?~������4�S�K�Te��Ib�������o1[�|:ox���/��Q�]��ʾT,����N��}������~7�U��ؓo���N��
1���~~�uL\J@e�������}/dr�'��b����������]��ޮp�_5����б�{���a|\���n�g��h��G��+��f�;S�3�grL�#��<�&P]?�?���y�����)V�ⷺ�q�|x���������2�С|�Rw�ϤS��Ej�N�?�S}�.7ڲBp��̦�Hr��?�^�	���Rjm�HBUeͶ��O��p7i.��A?���<���x���a߅���9ѓ��}�RS����W�G�:Y����J��&���0��%(�{i���Բ;��בrQ��d~���G�ү�Zat�!�4����dH�+Ԕb�>s�U���o-#Y]��{-�7�8	J]���I��F�[�1��6���l���Z���45�*X�^��9���F�"G��/��o�ѹ��f�3yBY�|���mMJ'x)�H�`f�ڿ��Tdsl0y��͉�߸��w4�F�蚉��͆?��uHb@^��e�Q ��W�5b�l��Pj��0�"���p�˗҃Y|rcϕ�4~Ue�: qDk��_MLT��UlQg�˼%u��~����lh�gs���K���^��/	�@�s�˘C����D���볥k}��	=��GH��ҪOU�$�T?��g3U�F��-[�l�ت5��vc��,�6b?�5��l�F��c�(֥=��ЦZس��;2�ˣK�{�<�S��*���쫍���x�
���-o���ENW�2���J���jI�^��Kϡɫ�����?�y7q8�%���B'1�,��M��%:��CU>C�=U1K^��j�<k(r�(p+����d5?ey�\d��Q��
kO��s3����q�|6��ٺqREk���zĕ��cj)�A�y6��[��n�1��#�o�=e�,���y�kf��`������!0�%l�|�};�p3y'bG��roD>�a )ʦh
�݅]���σQ�!���i:��p3U&z����}��4�+u��XuT4RV#|=����I ��[����l|�I,`z�T$�����*�q���ע{���bL�I��b��p�Hͭ���c+�^�b��X"X}���G�)<�����iI�L�.�3h17��c�ehR��������;6S�_���Y�M7�*{�#��������P����=M�87N͔[1�l���͍��fe�"G����fމ"��tQ�G���f܇ѩbsI�j��LȬ��ٝ��-k$�����d��e1�Vh=R����#M�o\�\�d���7��l{��&t��4���ury�x�r�ޮQ�T���Ǫu��4����Q��p�����X�1[�!�T�E0��_��F$hvk�k-𲀧�*��]MsOi������m��<�VZ�Y*Z�3ü&*�����b�jɦ�0dUQu5�#�)�{Y��/I���T�o2;9ޖio�����)w�W�]4{'����g�To;���|j�#Xe�Z�ؖ���Z#�M����r��֖kw	�U+n'��vw��=�J6O�Ƀ�wqXn��V�M'4e�\�9LO�
��ּZ<�1�[��N��st�⇒gJ��.&P@�j�=>J>�1W�~c�}j1��we
[�m\|f��B�-�߶�r��$��K�����^���x}��E�����2eP��F��z�r�0���^��d��N��{ޡ��5iS���W�jk�J0��6���T�~�r!�67k�Ko�C���~��@�ƴ��>��`Eb7`
9�aH�ܯ��:a�7:RC\��/��u����%멡�Pf��F������j��>U�h7��n�ݿ� h84��
.4F���c� ��cuI����]Z��V�n��靼wő�P����^�����;���T6M�n�E�x1��Y�S����{�!97�}�&d�Ƒ'S�*�#Q��X�:���2ļ)ɞ��O^� Uyf�`:N�Т]c��C�ՙiژ�7�p�UD*��M_����l:杤���#�"�_�#�o��F��7.��zU��
4ׯ�{�/Ja��TfX%��f��wG
��
��խ'N�g��7Om�o3�x�j�F���0�9��H+����9�}Up�{�� `�s��X�BT���5������3�Dq�Q�����v���8���c�p��������}����=������m��󪼸'JUc�qo�Y(���w)�3yœ̜f?����6��`��A�H�!I�4��j1��ؠ=P��g�+[O�$�3>eX6�ux�f��Y0�P� uZ���Z�,@u��['��)ļl���l��k׊o@�1�,�u���Ň(���WN���s<JnZIe(-�/���C�K,����S��Ν�����h��N?\v��s*{���m�uf]7+�{���!^R8]@���O�Bc(���������!�1�S(��^L��/s�?NK<�<�@��޷��q�'��Ƨ&LO��.�B�j�`������v�
^Jֳ�K����8��Ӣ^�|��F�r�	��80�+9�cN��q���.�-}Z����R0Ꝭvo��o��G�()3ʵ:uv	�����#Y��}�U�V��}�Tɲ4c���x2�n�'R}��5?�U<��X� 5��W���*�_-
w�ލ �Ǿ�{w����Z�y)VI�����*|� Yk��G��y����;m��"շ��t��e�^�^w2�Ui=�>ڞG����u+��U���6��2~���*�W�"�ni��ѱ�����	8�	N��������	M��G��W��±H�^��v�hsh��[^�M�ӗ_�8Jє+u��e����3 B���o;,��� ���V�O�����
�
.�ގ���-wL�=�qx�?���J����+��^V��H��/N�x){m���U�S�]�-u�u��=:��@��t���0����A���M#9�C(Z�ka����=��7��ڝ���S��˸��6i�}ƇZ0��%3olH|��58�Wz��䄥#sX��ͺkq0?ւ<.D5k����+�ā�7\�Bx���(fn����WN[W[y����n���%�!9$Yϻӿ�q�7pn3_�x�]��jlȵl��[�$��'��c74(1Gl���|j�U�mt'fzn�mf�?š5�q�������U���gU�ܭ����R�g���k�VQ�{�5[85�mX��}H�9G��TB9\)8�B�r �߹�S��;��o@�i�Ywg^�ƾ !-;!ޣ�Q�d�����
�fm��Y��_�sm	��K^�7��6�*#��U�6M�C��xu����Z�9'?v	"u��R��V�0(��25~�itUm;k?�|���2W"f���oP7���a����z��#�#8!�����L��ϊ�[�"�	7<j'M���"}Y�)0.�_'�O����z�5ea(.���l��R��V����9�J��g\Ay�|vl�u����.�ݯ�U�k"�C�{�,H��ߚrP�C�k��kl��2���ޛ�
>x\~-e\o�'�p�݄�>���*�y���]әh8�w4^U�&�p��S�H��m[I2�t>�lw6�t���uD��[����������:n3*���#X�ب�?W����R�������Y��f�˛�>��cu��cqt͛�����ԳC��s��x1-z�}*�P�K
U���4���i6�Ǻʄ�=���]C�%GAȱ�&)ȕ�<��� �i�T����@H��>5"]�	��[`)-�I�1>�	.$�̱Ǉ��C�ŭ�Mg2(O-'�O߬��6�d�N7Kj��;�YE���C,��_�E}���Hb��=`rF%����+�����nsL�:��N1����E����ً�q��I�[OԽ]tXm�O�RS7[�3���p�L�?+��;�&|�X!��fJf �U��ix��f�M��2���/�i#H�4�qA���"��&���d�{;Һ2d�b,�=WID��Ĉn��K�����)bxJ�+�9�e,�P!Ӵ��o��/����w��l�x�y��ӬXagو&_I��C47L��v|#.�,��ay5�;�hpK~.:�Ԗ�N,��u�-�QV�\+3Lq����a�:�ӆ����5T3\g�k��>��q���7��`�8^9`���*[�f����~Uکg�O�p���_G��sC�_M��<�E��,6�t/��=ߢꝿU�;1���z��)d:ڬO6_���3��G�W���5=�q�f-�Il���!�Yn�6�LХ��j�l�	i�4���i���X/]'|����Й��H�O��J�����+��ݏ�����%����zކ]�t_�&Ԇ���4IYW�B�].� p�t�@�7@��ʴрU/�A�-#�:���VoB�r&ZO���9x�����x��*��F��e��z��)NŠ7�<��r�@��m��.�g8n����z+5�^���̾�k�A}p�p� Iw��1����~��v<���*�7��<{��Eŋ��@�^n"�/-5r�Y�}Y���W�h3�3 L�"*�Fn����'�:��9H�u����Rbx�_�|�g�цm������/e�d7�:�F���^�6C�Y|P����M��䆁��>�����y�Bud��{�M��05TJ�4�dp�!po�����-�Pe`v��z���ۄ����0[��(�����R�(#A���r����cH���j���K<��l��GėR��:��Tᓣ)eoҡ6�9���I����[k&��^��x��U3����%��gQ����ns� �s��(�S�s/�����K��a���.���|�����G�z��RDN��:s/�!y8r�WW�0��б���n�1',�輺������/�+���Q���Ț�Ιqe��_]�;"�;�V�<@�� =.�QQ,��g�!�2�1�yu�[�+�|l���;?6�E��.��s|�.�
����!�A����'�d[�����|$��=��CH��\�	�����[���Jg��!y[O���٢�H��_7_�VC��i\�d�ԔWz�
�����d�|�r�3�y�FJwl�.��D�E�����h��l��h�S�B7�>L~h�[?ᷟ8̙��-�.���ۏ�D��e�uҧ����=���q��P �B��X�v����hn�5P
W����Z&Y��n|���n���^��R�e;�P5�c^��եB�g.!�=�
5�y��^���(�B�8��k�(^��_���D�g���Ck�͵le�W����ս��T͔ �iȉr���T	�Y|�=
4^��F��y�O�0m��b�oq �$�f��w�!��x�4��͵��mZzO;��gF��5�
V{�.�6��+�V�a����|���{ϑb����x鷱}\�w�y��ק<UY~�J�I{; �-&>:��cLv.~�+�����+E
�0ś��p����|"�k��%cjX��a�n����U�ӋQ�[��{˪%�z�}G6��A6�����;�]a�ٌ��)8���Щ���R+��3��~�i����������r���כ�����;4� �"s{F��<;T"ŋk������=�sU�g�Ha��	�a�=�i0��@?������V\�m3�mV@b�b��Z��أ�|�����g�����E��<�O+y���j.�vi�B_��r8ד�#��s�ԇ�
��6H�䏞����p�t>���` �(Z)����2�@!��yle�C����VϷu���ک;����1&_W�.E�p�/ae���3�Uu���bX�Yt�'���+�p�-˪�����1�L�Sp��zq�ucm~��9�0���uɄ���fH����/����`���7�s������.=�;'mi��Ƀ��5�H}��Dh֨�uY]������MMP�zޑj����طN]�Ң�D�K������i��t�����ks����|�]�N>�v�+��y�î�r�1.�!��P���� q����V��B-�
vvG�#��
�:p�f�M
쫄�����Z�?�LLS&�;�00`�w��8V(m��*"� �ʪ3
����q_-%�x$��G|~5��>&�o��d�Ad8Ya� 7:�)�����/u��N�{)�]��W7���Hf�`Jk�L��#����G��̜#��D���r������:��<���wy�L3�Ïv�g���ԝ�s���5��`�7VZ�
gu<ť��y��(��1�7��-�D��Ԥn}�<5����ob�7�$�k*b�����AYo�8bi�T$��v�m@����l~F�w:5A�.R���:JqP��$�v7F#\�9�l��H"zN[����$��}�DN��5a���^�p��{���+��}��?�آ`�A��*��{e:ϯ��f�ݥB}O�|+�1]�C��A�k�(�������ŗuf�t����q��%�ɢ�9,H��0�';�+���F碹@u?Hi�+���M"c�*{w��_�s�Iq�,uLWL�o.�H������}���D��W #���!��I�U����Q�1ý��9;�E�%�_�/�d�����
u))��;+ص>(ay��z`�WVV3F}�k����5A#?���j�"���?|x�C_RXh��P۰��ț�๛���ǚ_��cA1�����K��lWJB���u�˾�)�K����qN� xOÀ"�k�?��C`��7LK�&6�:oK�W���m�����6Ԁ�]՜�T�V�4e��k�)Q8���w|#F���o���f��n��>��O'bdԬ
�YƩ�������6�m���y��Nan�@Rm�*[��2c9��d�gUw�1�N:a�Ȃ<xn�č�9G���)�������˪���$Fw��ߘL�h�-�d����?�y�4>�Xz�f�>S`���z	z�C����Xv�3�M,?Ğf��k��~��g4ط)��ˌo�����-|1Q+��<�������Z#2�P���d?�})vY�fa7]o���n����1��E�y>|I(HCl�����k�0!��G%�h���^Q)�v��ۦ:�
�!���5��k�f{J�,�tr8���(W��H���f��>^u�y�����F��0 �9�2o �8��_V�]��g�*���M
8�.���\�ۯ88C��?�Qf����#�3K\�/B��44bc���7��-K��%G��Sg�ݲ�-�8mp;h��TӞ^�}���h��i�عu�(7��cn;m��Ѝ�y]��()k'��Ω�%$�,]�C�Ƶ��_��X]�?�3�)�+����mg1���a��KY?�����ɮNŮw���^-��<8�0�?�zu9�X����yo=_i6:Qw<��d�����4Y֣���������*��ܬ(�Xj
P�t#KG��A�	�-�`,
^IR��J���'�~u��4�R0���&��u`À���'2L�8k_���lʻU�Y����n:�v*Y�W�S�K�K<��7$o�(4���<z�XA�x������[�W�e���s+˚�P��Ǹ��kQ~QE���;e�=!�'��a��͓�ҡ��#��y��ja�ȑ׸�p����~��x��i~��{��ce��说��I�U6[E,c�󾶺� л�:y�洛cߋ&���d�.T4@B�Ȁ�Ы�{�kg�I	6�@/�n����$��1)ְ�P�����A-��%k�V#��LSg�139�ku��SR�*��w�.s��p������\�$2�ZU���~B��ɌQ�N>�	r�x�_��υ���=�*\�oO�S|~�@	_��^�P�߈̮��q�u�~A=�o�\�@'������wY�cOk�#����ꎐ9Qb�QZ>#V7�>��^�i?���HrT,_?ț�W��z`������\o��l�j�7ab��w�If����w��&����d��7Nji)�$%�u4�߷���N57�{�-���׋�z�2�x�D����45�J&�f>m5�Q,�K�;�b��_h��Ƹv����vU6��Ć�>���Ԫĥ�^�aS��G^�B����`����ʺKq�C+�e���o=4��6�/�2�_�U�=jӯ^�-�r޵�����0��ۖ �p����w'8�IqZ>�����o��)�Q����xcQT_��#��k���뎓{ݷ�6�tB���{���Vs\V�{�NV(cO&����5�	F0��	�i�7�I���~N:�J`��<�2�?���?��������^�n��te�F�[��:��<����e7�gS�S0�¤]#��t%wu*�}��M��,�Y8�ߜ�We���a[�a�ȃp̃Q���ͨ�1��w���됀�^�+L��Hl��5,Fb8�2Q��A[��_x|Պ�.ʔ�i�
0�UKH:����^�l:�=6���W4����t.텕ӮO|K�UF���3u��rp�ح2Pzͷ�5x��A����ubI��RR��!�TV��CCS�9}$}���	��*���>
��c�R5(8��% �h��Y�K�SNov�����҉y�n�X$erK���-"��.�1�n�8���=8�ߎR�m�(t���
���=�Dk�w���#F9\7�D�!Q�=?� �;�4� �b1�TfƱaQ�|J��~�ZN~Q���18�^C��a+
�E,��0�cI6��<b5a��z���t_>�^V�CwYݻ:~? �2�z�R̼L}��VL��liD���=��J�q7)�k���(�eЇ(���|�E�BȧC�.2��s�ï���.zqB���D��E�����U�mԠI�=}�,��Yfү��A׏D1��/^3����0���G�8��nr�~
N�H������LGǠU�N׮�'S�`Р���8k��Fk�X��f�Dú֣���ũ8�T���e�������nY���B���Tw63P��S�X:��X5(���Z*���-���(l�v��b���e�t��L2�6�?��{��7�9�9.q���׻���3��#98��7깅��|�S>�9*޳�&e��z�6jA�K&@O�^w0AT��IPA��S��^�����\c��w����
%�EE<E��b����ɫ*���gC3����uRuQ�e蘯ʬB�����r���Q�F<�G�\�B�,���w,R���gS�k�{�1��'c¡ڔIɡe�NB}� ��kS����F�"�vh����h%F�����Ļ�-��<E��*?���ґF�/�� �p`�8�<D1$Uq�@@��qz�LF/��J��� ��B�D��ܬ�R��{��@ςv�KƲ�J��03Sõ����4g��2���;���=���=�r�\-��;ւ������_�HE���7p#F9�mݩA�����{[h������6#_�;gP�.�G�o=�Z ~�a�{~Pc��I�r��<��"���jk�~u��Q#!�9l16ȣ��I���;�*���WqX|��v�n�j��Z�p�D>�Q6N�o�
XK/�`���Z	f||$g�tx�$�9��� z&d4 :�H}#����ǭ²���T���Y�~����ɠp�gE
�����ޛ��Sݳ�l�%wF��.������b�貚��u�oK�ϖ�D'�=z�������J��m#y�B/�6��Q�"�\���r\��70�OP��Ҭ6�X_��^�g���:�_q��s�_R�2�p'/�F�I�=���Ai�{�0�"0c�����bH��Y(�l�7�K9�t1��=h��	t;�;�«)��Fa��=���iF�cmT�QN����%~��m��/#��x�Y��眝�s �/��x������č�e���e7~�x�ܶ�~����-h�uqp��<;�R��|��6豓;�P/I*��n�[����{�g��_����r[Ͷ��~�Ty̯ሪ��9��r��깾
��0.N�9��7����q1#K�.�ت��ݓL4lR��} q�����[.�i|$��<������'X,�mu��'���c�4ru�2mTƄF���S��(�E��^���J��J��B!��`������Gπ��3�M-��)� ��m)���j"�g�^X�s��w����(Hb74����i��w�a���U��ԉf�<�
�E$��1�i�����]�t��6�ݛ�_�.�s�9�d&�w�=���а�\��2!�A0��o?c|g�ډhMɷ�~��7bD�}2H�v�tv�l��<1�d�f;�<a�	�R@��8o��|�|�S� ��˝�}�tQ}��/aZI���{�&�x��eUT��?�O"M���*ل@� �����;�|UڰbL�����|I��;Z���+ ��E���_�P�d���Ė�Ie}u�}ʩ�c<Ps1#�����PO����o���cp��i3������&�ā�C�vm������W���I�%$<�YQ)ö�y)�Z��8l�}�2�R�T�h�*cXQ�M�@cq�����x�*��
����$����e�frO�KP�p�{����r���P�B3E`e�~	���pP���<���/�I�U"�ܷf;��@ͅ�!�dƐE�Ҹַ]�6�u�޳��PfS�[�H�T��T§gʭ��E	2`�&kX����sAIo��!1 P��F!�+�d��J��xc��氯m��7 �d��M�}{:{@���oB�[XZ�Uƽ0̅�6<e�\9?� ��H=_�{ �_/E6���a�����i�ͷb5(S�����qQt�ۃ� �%
�� �JJ7�"�,)a"!)ݵ����HIw� K7,������~>���s��}]���!-�9Źq!֚��F���Q�y���i�Y�e�j��-����HhI�IPS�`�����6Ԕ�Xy�	ւYR�z���ɼ�<^����s�i�4�˦�#�fV�TS�@�<�W�&c�`M�@"%�t&&���`Zsǯ� F�NN��������+֫r�VO��(|P�&SJb�|j����B����w `�K�e]&{L��%��dD�������/bU ��8(W��vN� �\��W��r��U��M��?�64�3"j�^,x�m���II�T��@5_	�����Ë���9Q����h�\�z��l@�B��#�L1��\һ��/�X1�Ӕ������g�%�����"Rw�V]����	���� fI[���ج�È�w��Óא�ߪ�
�����i���sɧx7� c�-��6F3]YK�/�G�1n�K@M22HOX�)�%��N���Q�8���seD'Q��ڇ��U�`�ϰ�t�u��CO��ʫ���@��ʟ٣�C��UV��Ǹ�h&��"sF�S���o�)��K	8r!x6��8$�ڂd	�ͥ��k7�����Ɛ��g�4	�_��?��q�Y�ɳ�1:����kyB!R��P�=|���-~��ܻC̥��!0^M�H��v+�xաX��l�ZI�v$S7�;P(	�WA�'^���g�>��	�"K<ݤ$��Eo�Y`��uͲ��;q��'��8�ix�dW���O��=�$�u�����ń�Γz<� _�\\�sU�O�m� ~��X/����e��9{�]ѯ�CU�п�S�Yzt���o��7U�W��b{�,�%1_������dI��zP��_���·6�Pg
h,{w��·W�(�:�5LP����W�2��ۤz}K��B��'�xi�< �46�K�9�}����7�U��Fzŗ�<�7ƫ�	,S��u�g���9���{0��XA��u�ax����
��K	q`쓊�sgDWn�D3J�|4�����J�?��{����)oM��չ��Ե�$$μ��7��R������k���o"��a0�F!v'hK�n�� z­.=I��@��7d� ��&7���6��f0�8j19���v{cV�����J���o�9ʍ�m��Qa��g�h�s�X�S�.H&>!ǷnN�C!���̈́� �G���Ҩ]�q�8�˗���T��x���Qcum��]%��F�ü��ݢl؀DF�X��{�Q�\��m�6�!��Ө�aD�zLf��I�|�:-TbLf�K�Eh�pD ��(��h�l��� ���?w�b�1_�M���s�l0�lb����ߣ�{F7ΙQ�ǣ�=o����(+	�X!��n��G�z`m�r�i
0��aH�v%1�H��JȊ�˟I��- �����7��k^+�}�~��Z�����-s����%{�t�MlLI�ƹ��C�<.�d��P�?��=4�!Ubm!�X4H���Eא��Wn婉�/�
��B M�5������@���Q��:�,��$�s���xHH�V��w��k��ZI�f�@Cqݤ�`HDEY��h�U�~���Y�3rfEw��x�G�)�.]
����F�7D��|1��q@�&�(��jAI+��R��V�č�%C�3���ş�� PKU��	��3�*H���^[Х4�`�R����ȧ�:���~S�������|��2�������6�MQ�t̱v�r<�j�����N�04G��\�gf�&�����:���7 �y�eR/Z$/���L���j%M�1��4�cl���v�{���
��"uxs�����
��g� d��`Y��m[��7 �|�/�J�@]M��R��[k] K8/����OH4OiiY��aϿioO�9%,�M���y��Pkz���tY8�S%,3�}yF\���E�]r����|)'&�h�g��]V����v�Gq$�B� �h՘zp�:�&T��'�庯��4ӝ��l�܎����>����r�냥�r9OG&���[;���b�@h��r���6��7l�N|���z|�h�#$�.ԓ�F?쳸vvU�_K&�������_
�ye�$��X
�r�w!�p��3=-��
Y<�u��/> ����><g�F��A���>�O�sNCB��h5�7�A�ԲC0��"��3�+�q���|H
���ѽ��=I�ck�+��``F���+ r|Dv��\?��fd�����Z� (��fp��?F��k���>�'W�ƭ6�-�,���n	H����çUU^6���6ȝ`ǫ����8����֋�fR��!���R6MY���(�:ӝ�ֵI�-~�^�Ec(fN��c�W��{��)�<&��Y{���F7�s�-��0�4���m[���a��ĝ���9��)��2�Tn���>�Zs
(�T�������� [�A�j�%B� Y.�Ӓ��qa ��H��P��v�%_)�K:d#�A����}��j��)�-��3���_��Fʻl����8���`������w�I�U��Ψ�)~9� ��i�.����?T���P��ԃ�����`@�����N��T�s�"ϡ�ְv�yc�0�!Z�hX4qՀD���,&����i~d��5�̯w$���:��:�� nϵ������l��Z����%X��X��w�B���F�4+���s˒�ͅ5|����⯬|�����?�\���ֿP�{&����b��@n0O���g7� ��<�'6ɞ�� �Rg��P~o��Ng$H����Pk�K�h�0~�0�T��gҲ����弒����W<m�x�?�4➿��\ʑ�ؤ�ƫ���h�ǈ	d�$M3�=g8i8Dww+�-
�`�D1i�ʋ��c�)C�HO*��]�C�~��>��$�u�~[
��/䄐I/*:�6J�:��(k�d3��P�� ALxD7"68�s�x$-S
�U��ȃh��eU���Ld:���.�5S�J5�L�hQmyzL�5��~D~.���,�/�k���6%U�.���橨!�,�o[��8�8aec��i �3N#�7]O� ��F�9q�D�>��έ��	h�_j�z�H�:�^�E�$�G�\���)��߄[� ��-y^��O�R5��^�7Ib	���u���bZ��n�7�����)|��d$��](���Y�0x(���4Xc����Yp�
���cNd?���{���?E�?� o�j��~�9/����s��kU����B��q2�,�PzÃ�A����H(��P� o$���8��z�9��{W�Cx>n��d�P�$G���+���/n����Ȃjz��1\�%�ɛ�1l���q��7
Y�u��K��O �'��kK\�h�*���Au[^e�����򡋏�qTI60#���Q��&4�@��h�A���|�?F� h��%v�������q`ԋLd��\a&�e8EV��W���X��&�7�5��)*���a�bpo��b��S�>�a@�_1��&ʛ����Ow��`�ÿ�ͬ䉒��E+�����d�Vt��k�L�)KY�����K�7�
��h3��` �����fv���QkmXǙ$B�����0F���C�|}�^��~�oߚ#ܯv+����Җ�AnB|���L�L�*G����h�G�ַ�YZd_.W�dlԓ�?�'` A~�ʒ}��E
�H�B	N.�[ pN��U��,*3�������:;<�(�>��P��F��5�:@e(��Dv��N����m���6v�c�BI	��T���h��H��Fens��s����S<ؐ
��o�~���N��4���t�1VO
H˗o?|�D�vU|��q�:���c�%��5�1�l�7��~d��@��־�����k^�6���!>ѽ��e�z8�%w�!9b���R�� �����kÎ>�0A�>_��?�`G���7p�(��52u�$n�~�-n�]2
�ND�����̸�p���,Vq�>��bae���b)X25	!<p�
S3J�e	^%�������x�ziD�o��*�����x��y�OP	�=���6���>��C�4>��	~��j�I��/q��Ӟ5�g���ro��yVu�Vt\z�& ��c����u�r�����
�A�:ncg`)�Zr_m/����Ƚ�G�t���~H��X*m��o'�@㿉����~��m�z����A��<NQ�Z=}P�U�s���;S�k�шLq���P0|�z��s��Uh��P�ac~�_~Γл�ZY��P*�e� �\�>n� -�FP
{���Z5?X�7J*�Өf<EPB�_�(��@��`����TS�P��%�	H\$����h@����6�q�ă �ϡ���4��������O,4#߂�������A�b�z�A ��g�x �^8�8�돜y����ޝ/�B�r�'�oui&�P�觥�)�K����3�����kk���4nL�-��H#�L��&PǕ�F�P"\�ǅ,ZA�t�Ø���0Cm���c�N��ѫjSPہ�����;��U�ux�΃Y���-�.y�K|Gw �Bɨҙ�|E��v	L�R?�;h9Y-�b��v~:��#���^��u{�w��	Ȝ}�`�[�rp_��Ǟ��B;�'p/Y[ФG8��HT�I���_�v{��qeB�A��"t������D�.`!��l!jg�������j腎C�'����n�4�c��I���x�j�D ���lp/x[}R7���.z�֝������ʐUD���<k��>Ðp*%�����p��Bkr�ZO����7�^�ϳUO
��}[��i#;h�{�F��͇Z��0��}@�1��	�Z����H!������ ��"훓@V{���f�*�w���C�E��$&p/0�X@JY���9���Y�Sk^�_�,]ĮL4���jbՐ�5���Ӳ������í���Z�g��|� G}>ힼ9� ,�S��E���r �K�6�r윑�hD�`uˏڠ �`��R���oM�mC��m��fR��{h��1�A���p2��x���M�w>}@;u�{!6�8z&�{�gn�j�G�u_��^�����1ho ��k7H)��)�Q���<Y�m��QI �Y%��~ő1\�E#vڷM#n��
�'�mS�Z�v�j8а F�jh��f=�=�ƍvEV��ނȥP���K��ܵ^�+Q^mmn'g�N!�;��>��9��C�DQ�P0HPF�ê3��KM�m0�Zn�Dռ�hr|��)�8 �
6�b=�2b)y���R&�ò��ے���'>5���4�7R�o�JEq��2x8�b�-��r)F��n&��@��x`IdjF�v�9�$���d��Df47�q`�n�اhgvw�1�*d?�x��Zൠ�!'3{Ug�ě��ຕ[�3y��l����:fY��ц��Q^��_�'�:E&=�sF=$ގ�˅��0�gn;��0b�1$��<]ᒻ�&6h`�у��c���ב�C��k��U��?o�8bޢ��T�!��"=~�;����0� `�3P2��}G�
�)�gߢx �
�
�5t�t�����[�����_M����>��x��á��ò,�OG�3-�������5�𒾗}<�����ʹ�-q��ԃ�{�\��F�#I��]���0p�W:tn׃0����N��X c�W���z�g*pt! vg�y>�Q�v{1K?�hH���L0u������W�W.����r�Pm���vKtH�F�:L0L�"�ky�6���(�g*߁jٯ!�@Vz��P�֚�e�]�����V6��-�ЌȪỻ�%�r���:fAtޞ���%�*��B�cS��1p� +O��xq]��S���EUF1�h�^d�� ?��bm:�燹#}t~��Lr��[�}���򔰞'_�Y�y�	��*��f�B<&%X�t��*��'�#��Z,�� ��e/���}�����w��g(6��1��\˼P�(�Ĥ�٬ M�_Îf�2�Ə�oJ�|0�^�g�}�d�%k8��ih��p)��t?*T���C�U�{+��Z2s�	{�F2�ȶA��@e�7X[_��mB���m���M6�@B����:/$\�C�������]����la6e��X{��I	CM�����_����������ti�[�=�Cek���T��wx��w��l]�kS�{��#�\ ���h��^�Yt�`��%8�!���M��Rێ��R�ZS�����b�y�n���r�e���{���������iǶ�)��Ǻ@�m�[Ww��li�����mt�v����B�X���������aWQ�M�!qo�$w>�Z֯{ծ��Gz`0��` R^ğ��D�������6��c��Pl��;�l��j����TE�mJPS��W�-��Vy�Hm;�ؾ	�,��Wc��Ni[�aP������&%�\��^�꺻����vLץ�|R� ��$|�]���������$s�-&��#��Տ%��J���]��E�6@2]*oaS�l����Z7ASV՝e��m��~ɯ�r�j"ɨ������r��i��p<p��J�k9�k�F�_U��xņm)	
��pcC���}׷}�I����@���ı@0�c���;�]�$ʮ�"�S��Ed�Osɘ5�	�tf�櫛�ۃA��	m�����u�&,�6�ի����<Z�~/��~�D@�ژ!�k�)i;�7^�rWp%�S�މb-"�+������JN�?yΦ�Qc5�����j�y)����폓8����Ӆ�|D�Ӻ��Z� D��y,/l�86A�|o'^�.|�=��D]�JVW4�Y��إ՞}�N;��}!dY�0*>�8��ۺpwl�����du�Q�G�J �.��q�Q�ʙ�_��ٍ����a�Q �6�S�=�v���M(�k%z���:���:�|P}`�!ɩ���Y:
`�0�!��/��<.�ٿ[q*�����
�.��R���O�5^�ҿq�h�<}�y�-c�3A7s�Щ](
�X
,���`¼,v����RϴK�/�]}
�^�7�Ć�N�]/7:�f����s����=��]ʂ�@"�o�<>�_g�8������[�A�v��w ����J����&	+|�cR��F������Y�{/�A�z)��~6�'y�b���4�?Dq����}�r��5���c�+���u���_C�D�3x��0�6�����V������a���vM�4���q����g�_*l�ksJ$;%����
@ZY�o�jxR
�[�2F9V����k~ :0���(�E�������,"͕W$��^D��;��2S�7징�ƴ��T0j3��GV{Í����o�-�����(*�%�\i�%;e:>c���H����>�4���Y�J(y:��T%�k���l��I�8"H=�p_��3���WӾWx�fQͥ4�n^*vqY�`�]u�+7}���t�]+��9��b�Ҝl��0�Z��{E��~��'�J�{�:�{�P�8�i4��o'�t�˓�w���Ffw��Y
���������#�Q>�C�4�Kcb%`<�ґ t!�?�������6��P�'�s�' �f͕���
/Ӹ������2����.�u#^���ɴ����p�O�s�[vj4�o^pH�p��Ps>\���~!���:�=�7���o����,����3\wĊl]��+�&uzh��Z��� �P����k�عoG�օ u��^Ԙu���ZF��PR´�O{Z�b!2D�"�HD����ꉮ���~�벉)�ub��XN��׻N^�����3����翯bcb��ÄU�(E�ػA�W]����?�m�ΎW��sMM~�5l<����.��w���T-}^�N��I;%�x�FN"&���w�{q;i�Ck+�\9P���o��LƑl��a<O$=�A�G�Kf?Y7�N[s�VvYg���{}I�ȡ8������i��%;x��ktq����U$�@��qR5N4�_��0���Td+�=��ʪ���D#rH6�U���q�'ve)�Sl�tI���}�}]{��6aK�����2���Ogoqş�Or'[�T��
��b���G�}�o�!A��{��'=2��s��������kL�/hw'��N�3]G�s�̞�7<\�$eP�hr��;&��>r��^�.l��V��O{�+
Qtk"�� !��i�K�����=�w�$��5Z'rF���w���!�8Wĳ��u{�rq������oq���1��B���ڂFM�/*�(��)��㬢9�hr�)VgX��{�Z���ǰ�Z�����8��Q�9�1u����Mǃ.9�+���Z�YiZ�-HUA+�k��f^u�$��V��D�������﷋Mݦ��7)�3c?F'�/&����'+E*S!|�#S��ĽmL�����'�����]ы[��z�����!��\��ϥ���E&������1��e�~E�����ʨ�JYE��+����`�s��]�����ܼ�5?�M��"U��	"E����B57 �]2S$�������R�OKW)�|L����*O�O���{���z�}�Dfo�P��Z��ؠ��h�S���N�q�ˋ��ϒ���J�.�*�q�'2����9�U'�)R���Wgm]���PE�
��Y��k=�Ǻ'� �B��{1u�z�&:�ؖ*
�8���)\�z���[}����W>��h��M�ʦ��i9Y�ͅrm���OM|
�lk�W��ck#e,"|]��f>z�R�no�z{\��:�P�63�w��$�a�rN�c�{}f �GW��8- ��v&����
�_b���T��k�5�\�7GG��h*�'��X��Y��*`f�Y��搉��HW<�Wzz8px�^�Ơ#���:�k�6⁲!۸r��g�0��� ���cփC۷=��)���L�� ��Ϣ�-X՚�2燄%���A#���<�����6)CRk[�)���?Z�nN˚�E���憓p����d_��$ke�WK�������L��w}�Y�S���ʗ.�o'��I4=T*�)H3�#.R�(����9S5ߤfH0�7]�箧X��˧��Yp.B"�ܭ4��7�F0�O)Yz9��_ zr�{���������B������!"�x�K�k^��F��D����2>�~��ge�"�ە��浢��ւ^[�c=�X�U;3S����K;I�����V�
�K1LH/�})7�ہ:6�J��h� DH(�6s�i��;�>++k������1VUQyp�|�f�%{-s�X!�,�82g��:)�^����@�y�HHC�ߑ�zu��u�Ae{�胼`#�^t��YŨ$Ի
Ԩr��	U�����gc�?�\�F-AV�C��]�b�_��SfYJT-��d,���BA{�e�Rr��:8��X�4^Pޥ:&�[f��gy�6��YP�Ց9�w �ʱ�b�Z�/�@CϨ��l�բ�4^W���Zh�U^Tn���kՑK�%K��9�?K�j �v��o����kU?�Z����G�c�G]��UvEr�����ϟ 6z��&<�9��^�Xh���4��Ͻ���EA�f�ٔ���Y"7�DezV
��R�k�T�*y�U)��n��\�����-t��=���l�}�)Sja)�z���烆����G��)�3Qz�*�3l<����L�[As%`��8��R���?0$2��$!��:�N��j?�H�j�6D��l\������./��4������:��8��K���T�\��Z#�DpN=gÃ�G��S
��f�+��x�+���?�Z|�	H�5˦���q�wϛPR��)�M2�{	?|����{!�百e�Q5|;e�H
7����d��8'I���|��k�Q.$��g����S�?�0��5b3����P�>bjI���p�~��8�����9� ��n�[�zYsQ��S�	3��5�z�
��M�{��&�0�"�S�9Ę��D��PJ�.��"�# ���Q+t�y�/p#,R�26Ϊ�pe-s��_�>���zFD�0�9	ѝ���".nzCO8D �4j�aJ��ߞ۔�.�-M���N%3	R���я��+�Y�}c�sK:�)��Wŉ��I�z@��� ����a^Ǉ?�06�f���0��6nQ-<���g>���R^j�q��`p$��r�d��W񁍰W?�(�X�7^� ��kq�1�EGH�B��.z3�.�ŷ��ĳ���U��L�B]�;J3;4��@��pWXn\���O��wM@mV��B��4\h�ta�5�#�]���x/VkJwێ���rⰵF}!`JŨj|K$x5!j�m�kC־��x����"�X���h�焝]|��?�c�ٶknz� �~^�������k�c���U�y��ٷ�E↢&�+n+/���@H�8�E�f���,7m^��������Pڱ�1=�#{� �l��kk������U��Pl���N�YجU��d_z�U�n��C~���8�M�&ƺD�u�[E;x�o���\�EÎ���&o[��(���� Z�����H(�'4����:;��Cz�wl�F)�
�mڼ�xl=*[��d)e/Ta�7/V��+IՁYY�\�`5"0�ɟ�� ��+v��[)�k'':���oKg��#��6���k��M�)MuB�/�e�o}�bϥk>�c��Kc@m6x���<昜r�wݤ�U�g��݂q�@I-��6�����\�չ��Y�U�B��'�I��肑GU��oG]��c��K����M���y�6��{6������5��K xc�6ǋI�{����}b�C_m�][4lA�4nt2�y"�ٛ��Ȁ�cӕ�SV��Q���M��Gz�й��f�v�"tw��纱"0�@W؅S·��i��f��4��^���	ѵ�;D~a=��y�����Ŧ�d-��h�K�C�>[������U����zh�D8�"�1�i\��XM:�
a"rւ�AI\��c���-���1ƫC��k�s�=?��Q�S4k�Z�����k�'	���|iԨW�N{z~
�-q�9e����~9�$`�1|%� 4t��fڷ�N�ϟ�[eg����g��f�����e�Z��7�$���f�r[ts�m�����!D��	Ԥ�:��ڷȗ�B�	�H�ӥ����+���rK�L�i��tz�\�m��GQx���_�_�R����2�&�]~\L��]����_��6�`�VHE9|xK��5h�~pB�r0_� ޶].����p���Y~09��X-w|.�����>l�M��
NktR�b������uά�����WA�������Uћ�g����#�֗�mM��ra"�!Z?���)��Tʡj���<w�s4.7�i�dI�2��,�^3%p)�Y��E�G��Z��G�ᵤ����`O�BfJ�z��`���+ů�\�--R�R7?��p�����r�~@N��3S�W|vڎP4�/�]�.?.�Ӈ�R;�a�H��?�%9�������U`_���uʴ���6��BPF �x���c^�l����?�\�)ձn�0��gX���8��y�}�Zi@��>r��ō4��)�y���
e Gm,P.�b��¶���&Fxh"�,曽���35����P��7���J����W�~��R�E���Tu�n�y_���̟�xѱ�W-��v[��ܘ��s�GZH�p��C���ٚ�qW��I0��H���A��W#?��%l�
'��&딍X��ISZ�7�?�:#J���|�Fr���J����r/<�pѵ@��l�s��UͯM�Mt��Ԕ�O
��1n�-��ؔD���b��=^`%j�2��^�M[���.{��vmk'c!u�ꔤ��O�N7t^�
:(��b6#�1���**ۙx;���!p���V��.�|������B�e��j�u�M��2Vf��E�)u�d,v���w⺙-�V��;�p�^�rxDn8>>��
����akjG�m�?Q��}���o�����v��D����M�q]�%O.{y���u5_�3b�K�8D%�}%LT+�D��${K띃K}�&�%�W�L��BQ�N���XN�ח�̕�7p�뀠�j��Shm��%�����؍GεAӗQ���΍oM%����5��iJ�"P�I9+�\_p#�D''
M*��atj>�e�s�;[��!E�'�\8�L�[��+��R��_��
�F=�SU���:��t�W�7h�	�����bA�έվʯ6nt�k����>��5�TNC6d��O��Lm��|*�j�
�����/�iČd�'~��M�O�%l��Ew���wvnR	�F/N�<�%S�viKbc�}.�Dֹ�!y����8q��ݲ����`���jͻ�S拕*���#��}O� zC��>É!l"	X=�^C3��9���3�!K� �V)��}���=���8�Cf�K�غWm���Hɛ��� ���J@1g*����LU�МzjT��$�=Ev֞�U��H-�b=�,Ǜ�!�������go%a�:�ʧ�ş<͠WlR|�FO�����|$���*'n��#%�"����D��}L.*�L�v�݊��.v�c��O�����X��ݚ�y.CY��D!|���2/Q�˽|�[o�H�j��/M�[��&�Iu7�̯,N��+�;���3�̕L��U-�D	;��H��%������Ζ�E_=O಄ ��Pq>��e�<6A7���p�pas�y�-ݺRb�Ӂ����l#�m4�O���2ꈸ2�G��;^��o�q�aS�E�:XI�I�&��:�WEg���1o45�(QY����zLa���,5Ә�E0s�����A�7Xho�ܚ]�<��̇��Gv0;��.�]�8�':�8��=�a�_M&�-���_y����P�ss"�+��>�BI��0��V#\|˩GW����ja�q�EZ�U�㘔)��"���;zgq����:Z��X�X1GE'���N� �FEk�/SM#�$�G�߉:REy�'������a��Nb]�M���*]�:�jҡ�/�%����;F�61�x�VZI������,��L�,�iX�<N���V�s��f#�6�; P���T[����	�)H���x�"P�gS?a�y�ǭ���nr���u%8�W5K_�)��h�D�f�W��7��'%a����uG��1�W�T���8(���~�餋����
,^�濒c)��1�MAF��̓lxV�ă����.��J w�l�����Z{&�8?�ؓ��}�n-))�\��^��4~��
<�I:ߙ�'�n �bno9�6Y���˖��tcپ�-!ΌNvҿ5vSSP
�~檿�8�P�C*�tй�_���Ͷ�����/��X��EWQϣ��D�9���ŵV��=��Ro�߫�ZT��j'���ά��;������|j-���g5V�*�S���VR>�����4�J�<�m�g��%�[5ι���!�����_*�2�c���l^u��t�j:%����Z[�.<cƮV���Xݫ)�V���>t�fK���L9���S�J�#�EmL������T�o5�������<\;�����9.轁pUZ\/�������~i�\O[��T���2���	�����
�a�)�ƆZ{C(%L(\�~�G���Ĉ���ߧk�b5�Ν6Y�~��rG=������P��Pbt���G��[�v/�\}�q���{�mb����"��V	v�I�S��i"��x��I�-��	�`�G�v㦾���#���k���`�=�ٔ���#���[�f���������~lɶ~c,\��1�[�u�H�"���v�RH ��@�K��rܿ�� Xo�	̷F��v�>ipn.���y��u:�����?G���覵�3���2��I�� 
釂xCS#�]���l�io�	\x98�Sm��h"���S��^.�ۆ���dc�>�|b4� g#'�2���M�q:k_�о�XLeA�����uyW����+>5Ϻ�343m�����ov�nsv6���Q�1Y\�!l�>�X<O� �� �@��X[�-�&��Y�$�} b����`A�'�=P����������݈󆧍�9�E��iM��.Y�I|��}N"r
Awbp�=����;�������O�Os�T�֫_�f�&c��f��%=����	W�NC��k|&pb�Gb5m��%΂��N}����L}��-P�����O�_�1T���k�`8�l�egz�vz��Ru����뎎mf�k����3&螓q ������Y���&�Q%�J��i�cq6,�7A4�_��l�����O��V(�_� ty��71�`��ó/?���@Ʋ�����������sT���`B��H��{}���ʴ�sA���$�"	`m	F��?�Gz��ېj,^�!����Zn��l]�T����nV��G���|6���.�1�#=ui�=���S[-ec����h�2�G!}3�G϶kS�5s��Mw�	�r�=�(��ܖ��0�����╌��}=�WI(�_~��|�b�u�δC�5h��{^�R$5�K/��oՄ��������&č�8.�:4-1.4\�}���3��g����]L8f�L`=��P˄�3a�L��7>��+��ڝ.��M�߅������k�Bd�;���ż5�}�>�`���� ���M�!zq��ztX�!]wǩ*�x7�J��U%������~��sWO�M�f"#U��C��U�:��h�=\bذ[/�����|����{ff�>iZ>�s�UyW���?7/�3�/�7 *����n8�U[q�9��oZ}6�%ηQY�G����!������J��j� c�qPv���T	_�zF�
2X�^�c�Y�7ٰ�!R�(�N��΀��ٲo5���q��vCߎx=�YŶ��i�MB��ym����~�Q��n�ӕ�,�Q� _��eBWl����L[ݔ�]������6���b���wW�Z�
�J�K��:|��t:��J��+`\EN��[L]*���vA�]�Q���e�1X����y�1��l=���)�p!�7��SE��I;H���Ƣ�;�T�T�8a{�Б!�7�f�R�ʷ�a��%uСńm�����j��u�XO5ԩ1����68 g���Mg
~PB"��Z�̟��H�A�A�����T�̐+�r)(p����dϜb�j�l�����ݶ/�t�p�峬V��O� ���V�����B5<��X�5��Z�:�e(h�i�rI%� PǄ@z�od�����N/~��{���~Y�����ʲ#�%����zD�ӟ.v�=��U%�x��wߔ<����z�i��v�+�5�'�ۯ���l�Q���sI�����M��"�b� ��M���.Q޵�˳��w�u�W��=�0�:�_GjtSL���I�Y��SF|<�2�H��h`s'�Z|?]f��o�����X�̘ޗ�)���!�����"���b���]��X#�Kf~��Z/3�S~�G����b3�Si���~�p��$��i���O�j�}/s��Xt�C���ؕ]��|��ǗV/��ocP�7���Ik�*�xG��S;���9�,�H:6�t�O�*Vܿ��iWJ��)d������n�i+7(x����>����Ӳ�x�Ԡ��֨�)l����;".�7[�/��7%7�ۺ�y����<Yߪޅo���y�7Z&�c�}�CW>���h'c]��rź�RbdT��J���C��z��鶝�`���,�U�e�Tb7�Z���c� ��i@#(��f�ӏ�/f��S}u+F�$�����3���ː�w��~�Ǳ�ZN�[��o�7�EY���۾$-�PJ1X����q8��n����ka��C�4�H�d�o.2�Z�`R�_ˠ 1X�1��A��W��D�>�ue�`a��`m���e�xR���#�_�/l��xC�c��m�6��I��/������,D�	d����]���5�}�����i*�H��S>����4��B�z��^��q����~�ؔ�8<~����[φ<��iB���m�+�),sc�dLե����uQ�9�8�;�P�l���Ŝ!��~�t%�8�����%��^�<�Ϙ�z���!4Ҽk��-���D�x+�}����Д���9�"qY���9�@
��<U���>n��`�A��֨�~Fqn[[p�@��-����Q��nn�me>������g���_G��6#n�������r� )��Md����9827w7�@�}]�1S���	'G��e��BwX���Œq�]��e����%���0�V+�ǥ�4B��o��K��P�c�7�`ش�����3r��{�ߟ��������Yf��J���ħtl���0�P�v��7⾡��"���w�m`-���YYuD�7{�x͌0���g<�g?�"O�M�|��O��K�'@���S��yp��K6Q�^;r:��l��.���h�W�$朠�F.�b/����t�1}\Z5�
��Ð_&��fsRGzD���>�Ҽ��#�@.��u���v%�gI�ƛ�_ e�����R��ɢ]������r�I�y���B�e̟WU�i�Hl���\�����^noWU�,i�v��Iąi�1�WW�����T}��Qr!���׏�4B�N�Ib�֥��]fwB�NĽ/�������^R�	f���Yy�X��?|�O+S��1b��?��y���3}�~�]�6^<(Er+D���{h�J�KFJ�v~�v��W��� ��`�'��)4+��F>������"	�r�VV�j�S� ���u<��c�N��R~bb(4��.�X�gHj]�f�~��en��[۴��'sx�ç��-�h"�B�C��:��������4�A����]���kC��ǐ,F��u�aU�_� "H7@��n)�i�n%��;9t���[��A�����������3����k���Qn�n��������W� �<�K;��,��$h��еh�T,��Oሟ�2-�큯��-ꟹ}���nѨ�0����E��Tx��`D��-����r�C�6t�-�r�����-��m� �&u���u,�W��_0�bc�g�۫��9�=	f�6[�$-ILM����b�x#q���"悘f�rh��- �@לfúF���TL� ����%��ȃ����$���P7���ƖQ� �w%g_��y�݊~�*1�Pͻ���cf?I�~�U�z�"��|����Ƽ�G��~�����TOݬ�v�n�x�:"`���U�wR ��	�?��	�	���T0�� ��u�z���� �۞@ˏ��f�c�n��F���B�L�Fd�x��Wab��WO����L���G�u�g��>�Ir�[�,Q-!��I�6��BC�ݨJ������)���=Ꝣ:���X9��*Y���>��*�ʬ����X����e`��Ʒ���D_�ԟ�����,��� �~�����q�m)$<�&��~0�S�L�x�P��GKv�N�s���%F�}¼o ����pdy>W��!�k�?�ɰ�������~�-D��ӈ���t(]�+0pw`�zy;�d�{��������7��=�z�7��#��ʾ�O������ҕg(k�P��j�$`n��I�>�����{�;)W� �(�c5da;1���a��e-�,Lf�OC+	��no|J܁D�
1�+dF[�;]+���\G�HFsu���^G��&���-�&�z�rdh�=p�]���j�0�U��[�����k ��8�b�;�<��n�s��gٿ����������<M"��%��N6��?��v?v<�Xu�#ܡ��]���{��L>� �5}�T�pʵ�<����7��0z�)��l6�e��'���M,,>��i�$@Y.O ?~D��^� c{�K�ݛ����S7�7�/����K3�;�M�����Ht���'t�����aK/]�c�)r�����"�IfڱIC~s��ݠ�K�r����?�$�xR�5kOY�h�^�A�*����G������;ʭN�7*un9y��� ���$m���iQX� �������G��цS��Z
WA��������3�&~S%���6��O��� T�i{��>��I`Kk*��^�3C�B�lc�O�TE�=�ۤN�hGP��φ-꽓z�]�P�b���O#�3a~�Ԭ��8f�5K�j��2�\60��M�)(�;�D�5r �7� t�p'�0R�O��l=��x�n�;E'�'���'���������9` �Ϻ�1��L��j��֡P���'l��%h��$���I��Nk��~�Ӭ�͹� _&�=%g��!Z��n����4z�>C,.M��X#׳����D}Y1���<X|�"��6J-K�vA6Sy�Y(�����v��eo���HA躚��e)G(�L�.����LY�|zQ�;�v~=�=_��؜�ۡ@^;N�n���?�Q�����c}�X��J����r����_�O��g��3~&��HA��,b(˸�R��В�e<_��fzhz�GA�t˥�cCZ�G� U��iM���a`g�<sGr��0!~<��߀��M<C�=�����S��������0y��>�8��M���P����X�c\ ��y��D��,Ja�_vھ�n�j��1�fQ�_�o�$L��Xj�b�3Ѷz��^W_����Ir�&�t����O@�.	���x�c��̮�h�U�zr�<є�����}W��J�{��" W��$2�,�ҿ��)�H�����Ν��i��q��PP��pHmc~�CV�Cwn@K�#����ћҩ��B��N��t${��������ˮ���c|D�E�� ����4�x]�	������UӪ�d�~M����Yea���Y���"����ߪ����1��60�����(=5�=mN`6��$m!���ϭ��1N�9B�V2V죗��z�9��g
��ǧ�3�hl��ƴ☕�}�;L��#��xXiq�W�0��R�F?c)V�A=<R�C�2�v
;)����5MA`h�>�O��5��[������^�=>�X20jN�o[�R:��.����%l'zy��&���6|Ì�o}����@�} $���Qko��e����j�Nʯ�5M�*�
#���~"�<zk��݌	,����L���5K��<U0�2`t;M���Ҳ~�D 9��nD�o�g���t]���j1XKu
���N�/ݛ.����`;��ǖ�0o�c�_��o���L5Nl�d�L�\ !���!0�$i�NćY��?���Ȼ`-�a��%��t|�.����Q�x�O��m��>�a&���U��Y�40@���7�(��?��^G��m71[!乩�k'h���׮0H������%�`��rm3s��Sכ�W�p([t�	�ƵU�<�����TMm�=>�⹻�N�� ��|��6�.~И��Q�G����u�R:�~���=^�hX�U���R0U�p=�EK�_aX��|�A �yt��:p�|�Q�T�����@Gf{����<�:�q�և�b����[�2�CﳻR��FK�H_D��� �6�k�����k��Km$ v��R�I(ąϋNh6�ʱ3���_�9+��zxG%��/8�~|eS�<���*�  H�u(��!ˁF��b ]z2`�H�ȱ��81����3�-��=�;��9:�ߗ�$rt����۵�Q��q�˫&U �hU���)��+�PY�92�Ѫ\�{I�߅wH
��Ī=���% }�[w��}�*S����$V�8��
N�vu�m�C��9<�մ�TY97@�4�P���ּ�K/6�ּ��۴��(�Ċ��a��P�qV��E.'
�4�ږ�?�@%�{
l���	��k�rZ��D��9=��"@��+���W@��p ���)��߹�z@~/�tD��)�03��N��t��?���_���E���U�~��K�v��6���m�>p���;�Ѷ��[��H�'�2C��+n�⟔~5͢��p�/�u�������!�
��k������\I��8��y�I�!���Y�����/�W���`��%NW�`v����{��*�C~� U�ǚU�����wA��/��� i�j������5�����֯%9�*�&�|�S�a����΀�=M���w�A�~M��7i&�$�b3"�`{�����c`~�=���/D�~����
�X�R$��ơH���8�c=�Q�?��H���U53fOf"7o �4������f�U�4��YJ)��E�Ԏ�ݯ@�o>>5+����U<�:��������W���I·�������ം�w���8N;{6w@6(x�x���c=� e~DɈ#��X�73�k׏� �0�Hj�<�u��U�JG�9?�����{�;0�(5W�х�Ч%)��-�ߵ |5ͫ���'��O��q�Ӌ��>�?�1��l@�Ƽ �.� ���&�Љ���e%_μ���BfH������.��4��%�V	��J�)�w5g�,�4�T;d������O4 gMQ�.���Ȍ�N��5�<f�����{ó��>s�>�:n�Á�/Ȁ
c�T[�{Z�-�	 ��21R7�R�c�,+{�7z�3`h�.���h@�g&��o�7�4Ne:���RzMm*�E@d�C
�����i{~\�U����aa�2@�J�l�� �/Y?Ji���b�2X
6� я��/�(�M43:I���4m@�
��~8G��w��K�=;���Ӻ5�q��)����` P���7ˆ���[��F<��0u�w�P	���
�;'�V�L⦡��s��5V�&ǆ&�9��(@3�<궉qD���|A9�+�V�ɕ�w��Z��I=�����B9���ə_6R��\r�[gzU)3\�hz�����jg�Y���R޶ʁ��AE�A��;\]���x�n ��G|l�(V_fQt@V�z�ޢ	T�ez���_��l_�O�p�!�7���MB�6|=�S?&��R�q9�{�r��u�p�8����EL��h�+U�V�l��|� zRly��c�7\2��`��8U�/�����cϟ �/�=_��&!t����>Ia���V]rf�=X����b�s�l[�|�x��a!��^���p���N5P�?;O��ָ�����*?�iy-C3<CG"}g')m�����wQ����]\<��u��� �0�J�ϋ��I�lWR��º!mb踩sT�|>�LvW#�jB|��w߀9'��'�;�$_t����#j������DT��':���P����M��j�N�J�̂/�b��O���R��kP���?"$����ׄt�|w��{�쪵��I�h���v���_��v�#�5����o�-�oH��{NH�B�Z �()Z�d�(q��V��Fy2XU1_�3HOwO�
�҆q|��#Lމ�ta!q_��$3�T�N��}=���t��	psǄ��= P�Z1�7D ����n8�����G�;��K<`��}.����ӓ)�(���թ�~�I+�L��	�݌���/vE�~�AOF;�pEGBX�:����F�� �dO�=�>@����ٮq��.8�@Kj�3�B� s�mN�����I��RD)1�����0�FB�>�4	1���!�P�I���?�8�A*;��i��|ı٤�b��R_������L��e�iHc���rѸM?�g��H��*��r$���_a�l0�W�B�����8�丫$�����oY��Ot��`<�G��H&���p]�
��o���w�X?�g��R1D�D�Tdg�@=�,�9�p���k䬯~��������}�Х�B��죥�(��t�:ŭ�C��E��VM˻�:x:?j�X�&�;v�`��B_x�sa\���?����s)����G�(*��������s�.+������#4�œo��3��O�����CX<x�d��M�&�M��DmWHu,�a���M OG�앒$�d�u�\�,b6c�&�H;��#S?�Ep�v�c>{e�G��?�s�E8'�F�Oh���X�d�ѬbC2����#����>�j)��}e'�����"��n#IX���9"5�&��l��i���Op�R�0&6 {=8���؈�¨gDd�g�H���O�w��z�uhK4���?�u�T.g+�3ƃ�ƻY�g�eb��~{�N���"&s���p2B�	(��
~� ��~�����-���1��˒��������V*m�]2��C�7�Ρ4���ٵEZ�a���U���O�S�o��n�^_���96c�>��� 0'}�,�slW�U�4|�<K���޽��M?>��`�����©)R�EL %�L}�1�<@�j�0A<Q�Uڇd
����3�� ����LfJJ�X�;T�ނaw��w	w9�k_�w���q"�10څ;�ΔGx߷����]�����<=��)�M�������8x�j�I�Q���;_��~�CY]4HYP#8�k�EV�꺡�߼M��~c��k��{�<y Q����\���"z�t1�:�u�)�y��w����JA:�=	���f��>��f�?�8�5�o&��ږOR���tS}25����o!�M{�/F���R��޻6D����	�f�u_a3��˩H���� LʊR��w����R*~�ԝ\��yFi����A�Vp$���x�uD�"ߤ� �:�pPTuc���P���A#?ׅvQ\^�0�)%�-���(% �.Y'��\����`B|�l��㐱sz 1��_�OD�ǹ`X�/IG4Ғ�j �R�ɫ���j����&Omj��q-�<�XY�:!th5�T��O9FZ;���h_9�s��<������'���/��E�R�O7�.,u痘J��a��m 6u_"�pVuZOήѸ�E��sK����ބ�R<�5�7ࡃv��')xG|�,%��?F�h7����|�0!hQ��b��R��j�8�U���ߧ��m��{��1��g�+�$��{\3k�c 畫P\���""~g=�W���R{��Ud�����k������M��T����lB:��;?#�,��z�O&����Yfa}�\,k�D���*�m���FL[�(����5�l*��SLF:^���D��%����40�t�G����$�Wy��V���G�)9f�-!EGd��Y/'B��/WC���I��N!Q�|�}��������0��e�0�5ea���%*���Mi���J�tY����`��['��lF�|� `���(Ǆ�}�4 �:��ж�i7��=Q�������R��wv1ט���H�|�ҁ?͈�e/��mX�9�ڦ�x9�{��K@&�,�,��'��m�KO��4��5{ �(�',��˩�|j6\lVk�a�?,�;;G�P�S��/_ ��0qE*�b��Akx��g}���*���
Ӛ=p1~�g�@Y�z�]8\�6�i�/��Ã!fp��X��nώ� �i��!(��������Ys�4�iĿ%�/�z��g�t�[wb�I��?1R�k�d��Ab
�E�I'�D��ͅA��.d� ۲�C���O`�߶L���������r���F)	)=dh�F����d7o�r�Yʹw��aA���i�\H�QU�����%�������;��+5���^��g�
��7��K��ހ����()_X�K�#Xdoj��}]1
��YXy��2ā���(8��+�f#�NF�9K3!kg�
���oA-��`�����}�A��	��F�st��*��p�����:/x5ł�M�)%t�PJGO{?��9W�*p]L�юԘ[�����O��o��YV�젃@1�\J�U��,�dԒgTf��tJ?�悼����U!u��m�٧��������.��Y��T�C�B���G�f��v33���F�?5tHԓ��7�S��P�"��Np�rG35�`�&i-N�w~���y��J�BK��m�u��N/l�"6cE>^�1Ȃ�����X>�)HVA�G��e��:���,�75�&`����!��S��sr� l��x:|ʫJ����WD�V��$@�O��d��W�v?;o��Eڶ����2Ƽ
7h�#� #�c��"��� ��AJ���mX���K����ѥ�Q!팋pA�۵�%%Ԕ��RVH���=ղ�-�|�N�S-�-�+xx�H9���3{����س
;v�H��<tl��!��'�,.էFS v/�'�#��p;�n4�j������X�����%���|U-�� �����).+>���8�����t�>"��x���@�,���`�F 쌲�Ne�%���;�d�ibA_�/�0���O����oQO\((���v	��#���X�`��L��������e����;� LQe$6�Y>XO�ݯiD�As��xQ�aő�e���ؓ���M�A�wQmvz����*�#�iRԕ�Y'�G��M��F���o��Xmz:g�*�T���H��ֺ��wdE�.�X�v(����Y�ȼQS�]u�0qA�MCz���V�o	2��:k�p����M��F<E��@<�<O���,l���?�ԕ�иY� �V�#�ŭ[�Pl����`ZZ�,O\r��˕8MV��ޮ��6ёB�oRi98���9�}�{yO?�Sm^����@��W�����y���M��9�̖�V�0>iIN��Bv��'��Q���z�P�����
5z�"�?�}@9�u�s��d+�X�s�7Y�O,ĊϻłU��Z��SV)��#�vc�`!��.�*�`z#~�,k�~N	'%1�y�y�tJ\tV_��qZ����q:��ld`<����ǱJ�kSE���ɵa�a��wˏ/p��q�� G�=�?��p��!��-I����>��h��Of�Z��l��ܜxr��>�y�^��g\��1[�W��c��i�m�wP8L���׆ƹt��)�H�>  �������SL�Wk��E�=��H��L �%���Ը]��»�d��|-~���C0M�B������\>�S:�(������v��y�Q3A;��)�����$���ƀe>u5�<@�֔F�
`���|Cs�Ҕ��j�%�Q��c��e�'='�2k��+��1���e���:���1�"�� ���k�������dS��Z�f�n�y5�� fo�چ�ln�_���]��>�z^۫H1G�z�z��9L D1��2W�U���Q�|��]��(;�x����Cx|���1����SG(`�}�za���f�"V���E)��W�p[O����hr��jR&���H��)�Wjj�]�����G!äo{�;~+���
�B�N�@	f@�_uv}=�L*AJf��_aw��]E�0��������ļ�C:��+�P�SS2��>a�T0|�;Й)�s���de𛬔�>r���H�Ɨ��+C�d���`	@�ڝ�s�Ưt9'\6�ę�a>+��C$���wHo�����'�s@�M,���vV�����
f�����O����@|�U@QN�މZljh�n�+l�*�S��Nrjl�0���F� �ȝ
��No&��� Ǥ*����lV�m��a ��K��́Oy����޹[~���-��x����<lFD4��q��B���틣�G9
�Y�q)6V����}AB�Ч�28�l ��͹8
�74I����
V_}������P𪞫�2�7/�g@��ԏ�^��4*6���V��L��qp�R�'�J���TI�=��5wf~oon�i��������ne������7�T�g�-�(E�)��Ww�-�M,1�q�߷ӽD�U��m-�ҏ�ҏ�����|`:�HW�qrdU�P� �ff������H�]����F��n��x���a��]�"��5�-H�|����܃�J��27�)��9��We�EH��S�d 
���S�)hp�������O����s���S��h��p��f.Jcl���7�|0�"n��&��dM�O�=^��#Pp���66�lL��_�\�f8�$l&-o6+
%9E�x�!q�Y��,�ۓ�{�lD���r��ltw��Hw��.�	����?j�Ǚе�+�}\XH���i�C�t�!�B+tZ��?�0���T(����J�#;?�&����\e�����AFj�D���=��)H,�-
j���UR~e��t�6�J����8|<�tFo�]3Ézt9�;P���{`��XQ�WvR����!�
0���>w
<RR�P�ֵ
Dod¿�#>T6���q��c]���(������ͦ�g�ݎ��e]�ŚfO��XLz�ErES	��f"�#�~�����'@��3���:��%�/$�@yaU��[���;��w�����]bz��<�X�<����n'�k��%�Gv��G�T��ЛE��{w~>��$�@Z�.�0rE]��U�<����ݡ;�YD�|K�Y�ݦ�:ֽ2o� �"-��]�E�@k����Dn��"_}�^"ʶ2����J0Yg:���Յ�m��r�{|7qP�#v����ʗ�?�{����~Tp��b�b��RW�����.F�m},"��:����b���
N~�P��
m5 da��M/x�[wn1˦���G&�*hT a���5 ���4��'|��.ܬ~<���Us�eR!�Gc�Dur��%N[1ɀ�����W�e��u�b���{�#&���rƏ��#D ��� ��EQA���Ua�z�������1�4�l�۩��v��&��#Ne檭Pej�]��@��`��"�*��9*�0��w:K+����@TD�U�����y�p#�G�#���ĉ������$(bÍ����ThSMmB_�UO�9Wu��f�:�MN_My���G揑S��F3�Ǐ�����Ϲ;��i�ɠAf�Rk�9�kP��N&�L�����x�R�åF��vd��}ڹ+����?��x^��؏�ӡ��ް:"�:+1e=,�;��^����@�V��� 4��;����?�E(n��7�����k7	��:�ؠ+)w�^�b+��cT��
>T��9�Q���Ѧ�._A�'?�iQf�ی���p���>����2��G B�0�Q����#��#j�o�����4ړ
P��R�����B�4k=��]Zq�2��h�OP��(x �'~�%ޅ58�:��Mػ�����P�i1
'
i��*?�m�yc�V��p�e�f@~�\��e�/-��@l,����&4z%go�A�:���>\&<!"���P�� jmj�����Q�ȫ�~(�`װ�k�{@�Na`��Qߑ�:��J�%�z��  �G�Dk
"�m���ԇ{���v_p��5��1��d��4�d�@Y���M���m�ǩ	zc���$9P#�Cƴ$����Y�T�t����7�/@��'W�Λ�S`G�tK��.')ˋ<��'So�X�%.�NȀx��jǂ���H��F%���w.J|;�C�
��)n���s ���%K�aXA{6�aLB����i����b(3E�yz�)i�%�Pd��"��0����o5��)�]��P���hLɤ�]�@m�wye�b�hM
��F���V���9] E؄ ����u[J@7�lĴ'�a��z�s��;�7�%d�>��ϛ��$I��D�X\�8*)H	�1|i>J$_T�ٶ���fM�)��L�g�(BW����IB� �*�
��y\��  �7"7�lH���
��@�l(%�ڭW���`��	�ڟ��Ek��d�>ɯ4l[\���������j��f���^����ŁT�[MB5n���H&���:%��Л��G�L4��p�IU�����id��U�b�u� ����$e/�����7o���r���*+@�|��B.~.�c�8�9�F�$�Tf`8��MB��w�P�br]GY�H�g�Uk�_^�����^�(�C�ĥi��kFnYy�����_y8&��w���W��ع��<��F������xM��Oz���?�86�R�_'>���������2�/)!O
�	�'j<#��ۮ������<b1xY�S��*�fǝ0�+�R%���_U}�:A/�K|JC�ˉ8�mm̀��m&k�`����wadÖ��#N]c�~��y7�4�u��턃�EZ��J�̀qQ�.�@<�SF�˦;�h��S	(��dyo,�ྗZ	��9��4�A%g���i߸��j=�uD��`3��@"?c��}��vu�<J��Ԭ;ѷ]Z�>��i�s�C�^U��|�/�k���'�aߖ���R�t���R��ovo�/^m+��f�u��ja�Ɉ�wA���"(���\���'�~dŷ.��<�6䳿C�����$U�p�e>�w?'�=�V�����Ɇ��Z(}͋[�M���B^��R�x���ë���,������k)5��n�L���.>4q�.�G���b�����¤W��4ͯTҪ����5�I/K�����5e�w;��v��>+vI���E���UpPu�K0H�e~+��T�jGBG�����X{���	z��3	�؛B�0��AI� ZR�Sr���+B5���<)�ϸ�0�dTRN��5��捎�x9�n���W����f�4���k�f��=3EPFkU_�g��m�]�u�*7�I��S�t����GE�/�z�d�ob���3����%S��LS(D<7�"<VK1H|�׎�6�_�9`��uNk)g��><�@�X��ߔ�sE�_���Ӱp&�u�لZAd\�${�M�����i�#7����J�Z�g�= ��u�"<�[��������F�:������iȼ�͉Q�V������w�}t�4���z?�N��t����.}=}��f����>�F�7q���U���-��Y�멲��Ǖ���*�ǎ�Mk�+-ʡ��=��d������}�~j ZRj�;����;u����X(|�K��!Q�1��0-�L�{gBTH�b}８�\�����'�k��7�;�G�hT5w�Q������H��t����P]�h��P�n�/0o�뇭c�(l��;����o+��lV�V� ���>���n�qBxL_�Ff�ɉ4 �KFr�Lj'8O�W��]�՞���hK�y\E�.n"��2���m��^�����������D3<����rd1�|��_�c�<˫-v�UP�*�B��o��=�{%�����~�P��V�/�}�$F���;�<E�_�=Y#��������nm"�S������_�\����b����E�{��l���s�I��\Kr�`�2�uq*����ڂ Hk����u�	6�ڂ�ػ9��*���S�*x���9��R֮��xM��{I\��M�w���)��斪�磶l+Knq���"��XK���#�Sb>���6=�ɱ��B���u]�P��7m�Az2cb<���߷�H�Zy��SJRR�"��/���N/��4�>9C��5�˺@5��[�w_��l���仅������|o7�3(Ȣ�c['D��jb�e\0��ɯ<,�-2Ɗ��w������g�j�i�M����3{=���>ҡ�&z��Kv�h�F�҂<]kY$�UF�:|p�B<m��106�:e�z�����(�0�6�L7�F��n���S�{NL����X͑:�s���F�9�
u�|Пۙc��G�S�M=�>%8��Ļ��i�#��v�A��pV���r٢��ӄCڬ�٭l��b=��R��_Fճ�zvϢ�g��z��.�i�g�������Bh�m��{�G�D���%P$��8L���
w�S��g�˒F��{/�̙�]<h��ر��f�&�]5�oC�|�	ȥs9��VT�������q���������G|�z�m��8�������/r�ȝ]lZ��
�珉�'�~n�?�U��`ɕP�6��G3"A�T�/�~�1�V�`&�[�~�r>�
@����xD�v&�`��0�ąO��E\N�'�`gc�[�:$���F[Gwx�C3ԕkl�R��C���>z��������>�Վ�M�K���h#����2� �u���`�o���7�t�ʳ.��{�h�;��S��+I��Ѓ��e�����ܐ�g-Ȯ���B�},E��9.˸Re\�и��R��˼��T�}|�t���ӱ����㗙x(���
�U�p�(h��c\s���c�04K�:����<����Ւ�(~�7�=�>�r�B��[?ەB^\���?f-Էu�o��IP3�s�yU�.������[?gLt6�3$�������G�@7���<�f3��5���[~����z��	��J:�tU㇂�����Źz��Z���0�Cm�h�O	:RM/��2���_�A\>7լ��1I����g�u�>{˓��Ia�Ǥ��'eo>m�o]�)��y��br[k0J�?�g�\�A�8��][i�AJ�J��=ڟ�䆔�[3��8�C Ay��"��bF�(=G9����(>��;n݉��#��H3v��K���B9�P�N�;����d/o:j�Rw�xSYhĢ2���tl�nHcUX���݉���K�t'�Z����P:�2�w׈~�:^��8�/��&XE��Yc�-{���i��\ѣ���xS�g�$��͹��Y�4b#«�D�ݒ���J��5��٦���6I�����ȉ �N�������t�C��z4��w*ċq�#y=�ǜ�z/n{N� *��]��F�-YT�^�ˌ�qS���{�/�9ʋ�=�D�O^��V{��b(�PP[)^[����)����	(PE��H�`�v%T3��/N���o���	,�*����Ȓ���>zъ=1�J�\Y��e'30S��?��dƎ,~�" Z<t)�k^y�i�
0Wإ7�k��)����r����Sc�pl�WLs�.��j3��.?];ѽ<�Xle L_ݪ��4ȻSf#5B>/�&���X�I�]�R�a�ʜ�C����P��w�f@�^�?��BlY~�'���\�h��]��"��6���ʤ9|ns�Q��D��De�;�a����ؕe?����(�?��"rĆȜ�T�֭��m�sCIo�Ȫx;:�'��R�X���3"Wƚ�N�\I��UV)��kR��<� ����j���:���v:���S�L�������W��w��^�Ո��O{�/mM8-o����O\�	Q1$�Ë��шTqb�:�ٍ�N�8�Qac/{4���w��d-�A�2�h۝��UxT���2��N��}�+��Z���ZPM���%��j��$ҋ!�n���~;��%�Lak<K�򪓨%�ޝ�*n�b
�L�����NT��ȍ9�a���\��:&�l],a}qW����?�;ڷ	�����H'4�u�y�wt��/��Il�W&7�#�s�x��U��	���	�un �a/[��#]tJ�/��G#����!0�}k2�S��ͯzY	�&U�.X�Iuh!�i�+U��Z~��#��,�p�T5;y\i��|�<�}@N{|�
]�r?g��B=�r潌��!��P���鎭2��s;$'&�t[<Sa�U]�+R��cZ�-���6�h�8X	Ce���	����d���Sǉ/j�u�i-��s��tO�kH�i�Be�ߑ������,���;���ߧ`��5�iӖ좹�����pn����PHV�ҟ���!��S�RŔ)6pۅ��h���b�	�p��#"W��#!�d��\[��k�������	zz89����_/��,g�N�=.��R��R�¢�֏6�1���K�����С$k[j��N1���F�C����O�)�tJ&@�!�¡_+Q�&���j���f��f�<������:R�>�~a�P��o���T�Z�,��pwe=RoHW�U�Ђ�T����C�g���%&޻�o�$u�ds��Ea�)��4�0�.u��9ؗϖU�����1���W���gs$��X{�Wڇ'�+�>��y��W��-S�:�׵j�7���!�:_N�*�Z������YH�2���|4��r}O�i!���1�q�>E�^��c�hq�wڌ@������R�'���3ə	��p� ����ԉXa����7��b�vɓ�e�X����O�L坬�������f�!��H#8\�ULMTG�+�C!o�1-3�F-��H`�M�h��#y����4G����^E��2����e���G�50Nع��7�c�΢ӕ�\����M_�=�����N���7�c�D�m�+$��,(6�6�[z��w$���l���$J�7�{�+��q91��^�iV��k���ap?J{^���4�%g���Da"�;jͨ`dH���؁�G���G\��4٣Ȓ��Q�G�-/j�tf�%}��Ǧ>���x��O1{;ߙi�
��_/�C����ug�T���a�{�/�P�����������)]�2W��������C��%20L��bb/�/�2�p w�娿�3�e�*�R ,p8]HCۚa�l�xw�$b��!��=`�������1�o$A�D���*���IȚ����Z=t+˦�"���䗆�!�%-&��XѦ�agQ��}��Q���> <��� ��G-`se��l�B��օp�e@6T����h�Å ����2�[��2r#�#
�,mp�Z�t�O Aqe�"��c�s2&��>�[�������\�z���	��R��}�6��3��XN~�>޶��]oz.��p"�J�����V�n<�L��v�����Pk�V/�����Ҏ�z�E:�4�erC�8-�OJ�b��2x�/z�
Ͱ�Ŷ���g~�0�4�<I�;q�{2V�Dj�a�i_7	Q߾���b���ʲFޜ��\�F��R+j�@ A��W�)KM�<i���޵�d���duJ��V�̋�������<��m���s��\e�\R�tl�����QRR��k ?�r$Vyl�@e�:dd!���Oh?ͩI�g�8�s#�Er�A�&��S���+{S���8>�
9Q��1��+Z���x��������t��Q0�i!�����V��d�z�涴Ė��:��V�s/<��N����A?k}���:Y�y�zפyӯJ�9���'���Ӿ�K�nǑJQ��T����x�iQ�������*�	���Y�'����kC���Ƿo�T'ၶ���p�����!9��K�l�_�٫!�"����Ԥ`����&@/T��exq��oȭ�N=Hl� -S6���0�J٥�)[���%=�������8����S��+SLV�!��)��%!�VQ�!��6��5��sE#ǵ}��:ޙ���k������KJ8�v�3�v�
��׌��٫��lj�g�������-?+�[����J���˻�$~-�%��-���_����N�4��j�^�7����㾩�PEv/��+���O#�B?��v�4�17I��8G���D�mex�n"�4����[��������%�(��Z\�,����^�r}�&Mn��6>澯�8CO��:�
�n`��!�V�-*��|�0=�����y�s�?q�{���R���_��k�0T#ޅq�ƥ�|�$7�r,��`���_�sF�`T!��Ý��]ա�`Eٴn��a�u�1ػ;]����(����､-���z����|����R�X���7΄�lbyŏ��7��~e�s�D����H�p`�l_2�y��O�sݹs(l(@�h�v��a�%as>��3	v�f<�\oqA�ށW)oR|y�x���w�1�ьpcs!=5��G��4��
}����t�RN���Ҟ��s�����AZ�šV�%����I-Ӯ|�D�tl���ȭ�W�V�����"�G���T��w�����z�A���5�ʁ�h��TΟ
u<@ma<l\t���wO1����]X�󩋝꟩��i�8�!R�������?�2,��{{ i�n)A�n	E��:FDR���p���!d��;�3���_�_$�^{�uǚ�9���������.�鲹~:���ʪ�����/��ɠS�y8��R�g�%4�VN��5}��\`�S{3�(�8W����E���v�*9���E.V��;dv���)^g0j��R��:aG%����A�P���P�^��� �+?�+�e� ~�:g�� ���N�Q�;,d^���PvE�bW �]Q]����>P�n�E�I4�}����h�<���%�w���N���K�%|�"����pbW*�zB��@�u��ɐ}[j$���o�U彅����uSCtV���37�f���z�
rn<���g1�ȴj�=����D?C88�{\�G��ۀ:}'��>�s,�䁎Y��] )e�Y�V~7"���e���Ϫ	��L����^��p��-�HCh���u(s�	q��s������c���Z[v��.�]���w��P[��k��I[b]X���L�+A`�,s�{E�`˙�쩰`�9�w2�q��[2:�B�#�r�q?�6}^�^v�.E������oK���g����a�{�fJS��
�������=��|<?�-x�VAs����ճ�vGu�8&�2� 2vF2��U�@��;���X����|�J�ħK�z�����y5��3^���l��H�!),�h�E����1S�dH��.t]F�+ey�(ſ
r �6�9Lr�����Lt����s�I��;ě�h=o2ء�}�vW�_�3��~�������:*�x�J�.��?�O$�L�YM��.�;��\	���1�;/�9���i¢�k����	#ƊV47��D��/_���[l�n�AFs�x};ᬇ>����S��4�]X��i�u�|ѽC^^�kG��3r�/8T����=�Jγ��@2���3�D�A]�c�!˺�+zkB�ì�*|w����)R�M�*,��fO�+��V���&�+@+ˍ�
[xH� ��^��<�֞B
-��dU�[��w����ſrpV�����w�q�i�W�SF��~3^�H�l��QR�G�+d,����߿�8��/,�_B(ܮt�����7j��Z��a������{�M��.V�ُ�OS��%�V�*��+�g'!X��jk�>4�绂o)�،~q���H�AZ�aL�5�Jxf\�ט�t�	�J݀^|ы9�GP����ge�ɬ�<�8�yQN}1.)���OD�hd�Z�p�Ob�W�22̕(��,��P�ײ1-����|��:�A��t���1�paC�7�e�@�2�k�(	�W!�2f��ڰSY=�$��~f���-7��ظ�h�p���yq���%���H�E��j
ǒ$נ�Ǭ��$*z�y6H���_���M�їlu�Dm���p�IvZ�M���0�"D4	�K�xɈ������i�X����L]8�}��Ҋ��WOp蒅��0�R���ߔe�vp Z���^X͉�y{ǊDa\Pҷ�5�<��G�9��~O�A�
� �蔐fh�u�-`�Ȏ�ʹ�c�n-�۩&(��,����Q��C�ć�:G7=�k%#��<�W���Y[a��ơ
۶�vc Y}��[��[~�\W�m��Y���4W�}=�s��A�ar�'�G�|��DA��tө��2W葤�}Or��s�r�j�r��k�����0����>��r�v��:KYg�����L��uA"��=�3��F|���.Mi7,�t�tɫjm�N�f�b���qM]����#�Gr2z3�_�,Q�a�f��s��@Gn>���$7��:F@�܍�����l�o���N��|��a���'��ә���Yl���2sZoF�[t��P��Ք�<�c��
e��G|�x�/9`�n��P�a�70��5Z�Q'<wΏ�ns0����ĝ��>ƺy��M��涪~EH���+Ţ��Δ(��ֺ؂I�brLc�oq �\�Q|%��Ʈ�u������j���t�����MWֺ�p�����pCv�r�W�_�6�
�f�-�_`�����"^�z�������R�
o77-�B����[$*Z��';�0�'�%�9����ہS�l��jn���-]x_d���1w�V�]���������(�O���'�v����TH�{\T�9&�J��Ɲ񴼦�¿�/�0��_�ا�;^��C��.V���$w�_����t���`�~?�c�S9P�Ypì����cD���i\rEjZ�x+%�0g^�n۝]�Rfj`��FA�HW{2`c��i���A�A�vU�V�v?J�AZ�g���!(ԯ�y�p�D���MIi�p���}zu�W�ޒ	Ɩm��^��b6؈�GF������X�#����<��蛍݌�C_���u��G�,��~����ma�LjOr���t �=Ix�Z�� yM�p�KN��1 e^ګ�|�,1�g�dK�����z��6��_��Ҟ<��_H�G�V�����C\�������f*�?܍��b�0����/�(�\s�5�O��8pu�ՄF-���M_�J�h*�跟:�Lz��#�C��T��2���,�ء�UB|��5�_-���%���T�L��ڴ�|O��k�]c��ɑ��'&ny�EW�?m�H!O����:7��x�=0�:�������UI sN�3�M��,��oq%ԙ�W��h�T����G�E�-�Z�j�X��G���P"��~0+
��hP_����x��@=�+���������z�噆���<���؆p�����$+�����["�|�
1\�l��1*%dl4J4,�6#62��O�7f8]z�8 �#�	� �����G4ԏA�5������+D�Č^光�'���z�h������'z]hU��b���i��9c(ܭ�Ok�p�7�1�/B�8+�S�=�dK��X��+�J�⛘]�i|��IZuX>���2~��zi�^直S����ʽ����B60�#'ϣ5$�Ҡ��1���_N��E>��hY3��R�g��^��G�`K��ތ��
Q6	�!��?�ң��ٶpQ�vp�����B���Nګ���})͈�l�{��N�atp�۲"�K��}̶HY\){��C�MT��ηK�
�W�����*�
"A?�[��l{��F���Y����ؚ�%uf��݇xn���S"Y'z?l����jy Zm5����2#��P�ˊ������{HS 2�O�L�j2�"?�Y���œ�цd�@A[#*�स�6pb�����\�ֺ�,��)����j[���o��`tO�y=�q�{7�t�Y���=U=mq�����GTJ@�S�jڸ�����#��%��2 �N��������P�F%�}}�	���FQ&�����lC_Edc1)��B���^To;��K{ `6�b;6e�������Z�(w���x\���w;�`t��I�f�ala��`/p�l&>>-�����orD�����?��2r����<�Л�?:���uC1B�_Q�B�2��Ľ'�������RP��T��6
�Lb�Y"��%��m�sAX>Y4'� �>��H 	/�>	P����j���VWM���4������Ι�x�<�%�]��L=�
PB����pw��I�;:����'Э�v§G�&��W��$���"~�SVt�`�+{�%O���G����'&�eT��b��JoI(W\�ۇ�i�!�k��'lG?���W_[�Y8�}sR����X�o.�������b��*���/a_p&y�7i���~S�$�5��W���>{��S�`BI�'.D~~El�͂�j4Q�ǐy N{��T�Z��@�&����ݘ�M9����,ӡ!�)h���8L�&!Wǐ��eC߾�L����q�燖A��[�,�{2S���!_+�L��`��b�x�\�|Sv9s��N����l��2As
WW�	?J:b2]��<%{�ǰ&�����\ٿ��}�;3�l~���!r��GC�Ȼ[�W;8�����LaUb�Pi;a~�L���|l�r��Y`���lٍ3�w` �ŋ�\��r��N2���@ά
v\,F�OL+��li�R���*ʸ~a��
$�`f�Rq'����6=��g�Zy�qOwj�D�ſ���r��E�,�{;j��g7����k1o�6�T��P��y��O$&�����Ipo��2��ox�ZҀ*�Vӟ ����M���J�A����&3,u'	�� =���4��]�Dx g�}�.�[���͋�Z;���"":S�J��0{N,~��Һ�B�g�sd��'��UL%8���~��E���r���81��� Ij�<�����.�1�!���B���U0�r����r6k�3��֢*��O�d������l�Q2�v�ˉ�P�D���B4��n#ꑜ�QK#�Y�RH�/���x�b1u´�w���^�:jB(o�W3g�#20ɕ6�R�Ÿȩ��^�cЗ�o�c�,�|������5�l��{'�@�#�cd�Q����f�oVS:o��"�}/��PE6G��X��m��{k�FXEP��e�qSR�/�+��v0א��M��x��ߦ"��S�k��AԄ�$a��u/f�b;�2�vw�v��X����G+ݍ���Ɓ:-5HN��]�x� �TU6�Q#�H����e9�5ӷ:g�HB�e��f���F��Ԙ<��.bvE��z0�	U��>ge�����*����{@�ף��~��ss�c���EP���,�X�\ɳ__���+���@%��_��]���p�?���U@F�K��k�G"���kN�f�K�I����l���m�&#���q`,�_.����>Q�	/����A�*��/�m���Q�o��/,�W#=���0�Ob8�eX�k��iW�R�"n����$�i��Np��F�?>�`��6���(0�b��c����#k�0i�E�X���j�^�;D��6�Kc����]IC9����w��r� ���~"�k�V���K-�N
U�	¨�?	Ș,T@`GFiV=	Hc@�c_vM�:�a9!:4>�<-���� gE]�Л.���^ԓ`kf
iS�]j���d��00��&�N�	:L�?*h��(j�5_��	�5 9���n>1�=}�M�B�8�s�!ѫ$�k�[�*%���*���&�� ��c�~ŧ�i1z��]4����N$#+b�`e~�Ú�v]�WK'��ɲ�N�.�͂���G��$<Y�1g
c���V
�ԭ;�H뙙�F�I>˒i��5{���߅	p�L����|S(�����`�.=��
�܈A���Y�\���$Z�۴������ތO��s���A�9=8�~��D)Nbhby����B�w:fA�O=ċ>c��B��������W4ͯ����1�������hg�;8���M�1=�n���.���~�����4;�m���Zm�(����;a��Y��O�X���[Ѱ<�V#J�a�P�J�㮋��JfA��c�}S��g߮u�g����Wi��'�+9�=R���i�x�T��F�ӹ�e��8~fW�ҳT��� -��J����2��O`�M�h�[��α���KO$�hԁ�Jc��0��5�w�������ރ�Ɉ�t���v��	�mU�'����c���{�@����%ѫ�jm���"a�%׍�LDA�,��v�K
 M�U4�Q!�\��¦��e@c�ʸ�o���w��͡������/�y^I��b�s3����`5*|�.𙛴����=7���&���l*�����4���� �$����Ƞ�8p��yU-NF �_�,�@P��١Aƶ���(@"��'v5�C��B�����R+�^��eF�M�o:���Œ
�F�g�=�d"#��1�)^L�@��3���������t�,��l��HŒ��5�B�na�?ї$��ser�G���_�~�k-Y��`�0�QQ?{N���n("���$;|��C���u�B9�;� �
�PW�����S�Oaw18�-͏��]|�����k9*J_�J`�T�b�yo �|�F��{55ܼj��K\�|�{�I��6l���
��bX��P��o"�}OY��Z���q�T
<kR|��Bɩ���!�Y
	��z��9��RW���(��X'uVKys���z?�fH��zy�����,�����e�ël�l6�B�����$�g�C+m�[�k=����(�s�����G������wo�*n���g�;878k��
�g��w���o7L,��	�[fF��N<A!n+�OS֪a��rd8���}�8���~-vzwD!����Wc�6N�'�T�;�W�-����9,Mw�Ӵ��Qb;�N;*l@.+Ș|<��oS����Ŵ��h����=X��,HC��SG"c>����K=*rЩH=������[�Έ��;�4�V<� !�!����:6p4�ԨGx�*ж�]����dH,������s[X%��E�q�D4�i�{s�W5����$B�;Gۘ	&��@�LqB��i�DI�;����ۜW��P�4�8�]�[�b��}x��W�k�Ku���S��:x��/q/e>�1��1utC��E��O+l���~�1BM.7Ud�$� ��4j�w�&���p�lÊ3�R����r9EL�P4hiD1U�X3;垺M.�;:
��`?��c���K�4ش�IQ�, 	�|\K��>A�+@5���3���m�SQ$�"ϯ�fC�
��(/(5�睺r�lT���_!��́�=�_�!+i���W�<��9�6%p��-*��ʍ��F4���W^EU����HU���j��'�B4�lpM�����-�����F��[�(e�[VE��:X��9����h�%T[s!�]���9bB#@�Z[G�9\��cEȷ �\RGKԚ����޺�}*��G/���D���أ��1�w9�����_k����
�7�Y��7kP�B���ȽJ�|�$���]ߋ4uuK8z�~D���92)C�u�޺[p�"���1�+����Ά�$�>8TO.�{e3q*.|�����"{�w�����=	CK�"�)�G-�g�j�9 �R�&nF�T�
ʾʡb�Y��܁�A*��`*ǀi���.�t�u|����q��7��/����&6�� S/��N8��}�f���;�I��=a��"�F0��,اX/��HY���쫆1Gq�OCi�� A0���_�������n��	S�����D\<��t,}m�����𺭾�d:X�=
0	��Ś�6�h�Y@`�tYMC���$�"��i�M���/"}�(C���R���bȺ/�;y_��F�k.��7�v�2�oK�4?��zL�6gS,�4�=w�}$�@R�0]�2����OwGF RN��M2t�v$m*�E��y�k����
O��e�?����q&Be�3nf@�GK0�̈́�iG��`cz��؟ ��/rɭ�a��\���������r��"��A���/y1�>�崅&˂7`U4��M�s�s��u���Zڢ���4������q��޿�Q�:R�����`x�A�����c���䯛w/^yh0�z� ��ehd̋��74��$[�IjX�a���S.�t5�>�~
��	ܵN���1����^����̑�ۨ�&����Hc$�NJ�V`G�51���(*˛WA|7J�����=�G�B� ��Y�ѵ�Q�z��h�+f�r&���}��{v��5�>i�:���&���]���%F��Br�ɺ��Òa��'�'t����fs[F;d�HC��U����Xb茥�)z�!}H����;~E�Nz,Ж ���Z�#�_���pA��/�aO$�"UPm;����S�is�t���Mf����̄�3O~��votĢ�G�M�Z3�𻟾 D� �Ԍ�~�h���7EVw+�P�L��X^�Ѳ�����H��0R����{xP����X	9����pMPrC3��[U��׺9��F'!/{T7"�iam����Ź9>^�ϛ�0T�+oC��?t��s��Ō>�14M~+��'Ҝ*���ƀ1���+DU�․�_7Ph2��$@b���������)PGvJzd���ű"���zG�0N'�;�<ک�-��.t�&q�	I];N�J�{����yi%��tT�z���6�w"�O�N��.�����ֲ.W��� s�?)1N�^� v&��Z�Q�ŔwC�f�g07#ּ�)���ڝ����^��~���o���ħ��u�W��kz���g�����:�zt	s9{�t�-F��&m��N	��[�|9����4|M�EA�h�*�;��
�l�m�-+@6sgR�0��W�\p'9i-����s;z[)�����G���_�/�lun���㲽�bq�N�0��q�XQU��i�n�jgݾ��j����[ �j3�F=���O'���Pb=2��>�[�/�w��%�z�LAH|�9B}&�$�,y��p;,I�u��@1��Y�-�q�O_z�V:*��^c=]U�fLc+�\z��/J ��VϢ/��j��Rnۿʑ���_�7��>Cr����φ���GS��4ɖ�`!Ń�3��6���1X�Ӌ�D��A������W{�to���Yz)ʞ{"8����"ZxLO@�U��LS��Q}�8g���>��`�/�m�Yꪾ�*���k��)����7'6�A����tT��;sHc�J՝��%0�Ⱥ��x��^�S���R\<�̻0���>�G������Nv�ʦ,�;�b�b�}(������P�:�b-s�0�l��豁K��f�n!JCn����_��@�mN;�Yj�}���y^�TLf,CZ����+x�큨��*i�P�~�/�F�)���?�������J~�r�Yd�����>�
RfД��a���mq�s����YlDg�?���%�XI�l $�hcK�����������J"oV�oZ�̊���1��pX	 �C%�;?]��g�l�!4�j2%�^�\=F��U�ثq�QF��(Z�rKS��(�Բs����H����ו���:�/_�o�Q� �6�[����f��y��w�z0*���M# �AI�5"W6n������&GW��rp�f��w�c��~�00*�R�b�xI�>Y�����K�YN�7��zސ��>�2/]�3c��_���w��)��	��>Xg�t8��	1U��}��眨��-7�9$F*A"Y���Uߦ65 c5nB|M�稞hh0�w~۳���#:�H�����Z?�U�uLD.H�"�!y�ۘ�K�r�qy�>�c�?��o�а���_��\�1��& ]j��ڜ��=$4�E�?_��)�J��j|��Oc��k��ꇿ�w/��Y����V�iZSyL����V������A6�OL�ꭓ1�=o�\�uQ/��Vﮊc7Tz��ڒ�
�5��Hi��6�A���Q��X|"g6�sׅ�0�=�P$'��+��|�8�W���~.�I��O���Z���۳��(�g�K"��qL��v�ۻ��dV��4���G������1��Y�2*E����I��3Z�J�������#!���R�l(��6D�k�<��d��\�z� ��'[�Bw�����H�����dCP[3�<�,M�D�ǧ1թ��ʅ�Vy�q[�il5:)&�aL$�J�*PM~�j�l��Է�� 7%�����?Պ	��r�ucܣ���a���U�L/�yF�X���.�y��MA1��K^���$���s��=y�<�!�SNyG��5+`:fr�����	�oU+�-\.�\��z��A�|_B�����r�w��<#ƫǌ��Z��lY��?|�b��.,5�!�7�kU��`ɑbk���0k?cD�m�,3����b���E�^�H�`/^����%Nz?�ߜ��T�m�Q�ܫ"q8�o�b.-�D��n)������0�f�!���}2%�zN���G����h�z,rU�N�b�T�� ��<��8�7y-����Bd�+�9�����˾n��X��i�*��̄�
������3?�!�Kv������J�H���>E�,Ϯ�􅽈�=�I�u�'��:�q6�xl-�):�̷ͪ�Tq�?��6C<u5��1*5ԝ�6�@9�8p�6�hy�����'Q�7¢�l��-6q�N]�Oڅ"B-��z	�Z�s���Ƶ+N�ĩ�ĸK�0��M�j�f@"�*� �޲��2�F��rE�%�U����Py�I���s`�߹��[�� t�����΃�ɧA~䍹�S����2��F ��g��ЖJ�M�s#u��(���������r�`<Tɥ��'k��u{!��e�� �Z�g�{,��m�\G�s��,K�D���Ɛ�߀��{�����G�i$@`^��1�ѷ͚�Y���i� �9}P�@�Q�1��	�a��D�1����e�/��1mRޟ%��Tܕ/ ce/k��4HļsՀv��_�lE�eM�M��u~W,��t/��?���9o0���tf��;g/
�,���g3���:,�
{k�3�3�J��;����(3X'$y+��i"�����$+ܻ'�+���dW�A�M�� p��뿻kY/��g$C����尣�� �<gj���U��4���f�Dr�������� >��������đ������.���u��/4
�eh��/��~~{~H��C�q|�W	ϰ�����!D�,�������s�_�X1����!LZM+�]	`P(2ܟzMV�R)q�ZU+�������ɦc����P��,��L�5�f�m�.&K۱[����;}������׳h��X�)��>E}[f$�"Le��T����ɾaR�zQ�Z�!�8�� ��Ğ��V|5��=9}���ztn�;v=�������B!��zP��v+f��I�$���K���{�fx��yD�>;\�n�!�F��������0��p$�*�CV��bVN�/3~L��r�S��5� Io�e�g�Nꣷ�q`������\��nWj��e������H�m.����=R��k�y"��SE֩YD���anhF�㳄Ԟ~�C�q�0�R���*���w�:�3�NƋ�����*A��
�*sN�\�N�-��^�'��GIK-s�S��~kN�V�R����'&����lF�Xirˉ;�54�٤>�mv</�h�䕠s�����΁K�,�8#���-b�"`3��e����-9�<��[��w^Ç��3��|���Vx��`�+	m���BN��/UGzz���U =����D����J�|���x����m�ݏB��a���/}�)����u�7�j�@}�����hv^?�+�'*��Z�ڊ�m���'-�Z0�r��c׆u�;��,7"a4<e� /M�������g�K��Bi@��[��o�
4��l#�+��%k��Zr>�O�T��"ţ��_5do�q'�6a_�"�+�A��>G�R��5��֋3r��*	�Q���b9|eŖ7{�)��pt���Bi� �>�P0 ��������=�ҡ[�<n1�"D�E2?�񖰦�L�Q���XG����B�1xȕ21���'�c��\���-�?S�x��#j�f����ѿQ�`�]��EC�?��OA+Q�٘���.}�4;�����	�<$|���秃��T]f1�%�ǧ��?�7�`��D�\���	x��ؐ�J�,��}ɷ�u_B�N�@���ϧDG�Q�&�P�L��r���f�6�sɈ�ߢPI���b_oz�"J��5�l&������**t��g��a��M�Z�[B�b󒒜�:���m�0�J�1|c4JZ�j>��Z<oIzA��u��o3O6�q�?�����즭L��L\��ٌk��Ps5��}��ߡ�c�|KN�\¯+w���C�z��B�� z�_���񚀧����%?�g�k̓�>7��S�兏V�56�qS���L۴����K9J�;�:�Z�����++�uZ�Jث Y�Yw��X�L+i@��,񃘟����KO1(s�<[�^�IZ�>V���@S|2���ؿ��{��exY�f~�&eұ0X�����~��j=/ͫ-�����G�'���I6�'vl$	��=�߽Pa�SB��(u�6���䆝Ki)s������u�5R_Nj�'{�E��]�B��!�W��Χ%%l)�x�׳a�f��->�B������ƬKSvV��� e{
�7¼A?lH�KJKb��8䶸����߿�4_4�!˝eNr|�|�3n	G�
��R�AC�@<���㌰�Ȫӊ����Ds���a�Ǣ-={��`����H�^���ͱ���_�V�-�GS��E涼h�ޣI<k,Os0	�4�
�7Խ���<�J"�4���˻z�`cA,<l���f�'�am���ّu���=�rQ��n{��ZI�أ�]"o4�~Nb?+�u�
,Bx�N�0zhd���&�]u��"��el�-�^䯱!4���V2n�K���g�d�t�k���ӿ��P��fJ|��\��U��4~o�����tYń��+d��w�R�D����[�)͡]]�n�Oa�Φ����c�g��Qɀ��'=P}|�'i.�Nˆ���(��@�g~t?���7&��h�j���68.�b�N/ݳ�?�aJ����L�KSqJ�~����\<3�#�\����l ����綘㹃�m����O�R�����5!��gVo �q�O �A��X��F�&��Y~��j�Kf�al�`�Dg�a?�_I �u���$����ƻ[�ձJcH����K^�l����^��Bv�<�f}��n�>->�:������Y���7Z��?_���Z�#��~T�b�P��]�%�����4 (���,�)G��x��<��k μ�ǀ#���)��"�&0+��~9 Hg�9����8���x��2��Q�Z|3�m1z�{�R�ّ`�X1���9o5������ñ���#�<�N^n*�W:�.�����ǵO���^|���'H�E`6Yۂk��g
�~���U|����'" �oOTBC(�S���0�Q.^�8�-gM��"����/���kݮ-�q����s�����^�@�7�l-$�����Z#ՙ����W��g�Wa����Q5�Ԝ8#�+
��GP�yL]h��F>0�(R\v��^�ݷ{�D�Ot�8E�dK
zy�x���go��œ(u��EY${y�\�L|/���u������3c�9<N�x�X��Ӿ����O��d;V��%]_��|�u���D����'�,�޵$���3�5�ė�K6�;VYwc_\��ta�'
0�h����(�S2/���=�}����ѾR��ì��d�/'�ЁQY�1���}��%:�&�qs	r����	4�G'���^��`��RX�԰�ܲ�*�䱃N���W�DYGN��(������@���K���~|����O�iɅ �i��i��i��,��;R���Q"޿�w�#��}���;fޫ&�[��lZ���O�'����e�nA~�v�b��/�8�Ǣ�Ðw�CZ����1t�*S�e�jy�_����b�͒�-��O�rA�'�O��Se_�.1��~c7�R��:�70������G.�����W�~��@(�क़���
蚸I��Hp�ѳV���L���ԙ�����J�x�z!}α��͎�s��Zz�1����]��a�Q�d����������P���#]��N��^����^����I$�N{�[��������b��48��TW�yI������'����-�y-� �d��MG���P���X�Nw�.��w# ��f��Ƿ�{������,|ݦ�=Y����-WD�"RC��h$~ꪙ�����58`+�a,�E����I�i+�E�^<��6�E2�ᒑ����|��O�lz���W����(S8scb�3�'V�ڼ���NjtN��'�4ɪ�ܶu�y�}�e-2� I\T�KT�9&2��8P���T }޽�Eem5�B��AS��F�)!G�e[q�I�T�E�kX����mm~X�뢉Mb=s��=1�I�4g߽bz�����t�����.�f�}�
���X��4g2��;G���N����v�U�k8�u�W�zE���O-O�C4Cqv�C��b�C�'H�D,~�v;��� *Iѳ���q�ؘ'�k���93*�P�b��&��W I���t�nG���6�1�<��0�il���&�G0b|��)�u ��Q����������.�T�E���tD{ݼ�$��"�,���^�68oH�ڢH.G�_CC
��`��+{#9r��eސ或o�F�[.��q��V�JXZud��>q����#{�L�T`Fy��+�^�[0�WRF��;E+a��s@�Yc���@_ҽ�f �>Ћ� ڛ����Ԯz�8D3���:�-��3jmR�L���7�S��?3��ؤw�}��iMI��Ii�zǨo�6��/� �x��<����D�7�k6��@A[mT��̆v�[���sR�V���W�BIE�fR2��K�����>O&�{�u�[:��<�`��ŁA}�����1� gՠ �ջt�����7�K�G��%*�SM�~1��P5���[8�d����n �5q�;@L�L�P\ƩZK �I�i�K�8i�;�Lww�H��:��s�������Z'�w�͞f("w�e ����{ ��ؼ:ۮ��\Lh�����MYn�hx�K�u�W��e�8βϓ9�ځ��?u��o���l�Wǌ��:|)`����Ҵ}�:]�]ܸ*�+T��TV�K��e�C��r5�<-�x����e�P�g�x��w�U�w�[�jk��1�����o�XnÚo	M/��E���%x`T��C�o�=�mQ��ʃg�(��RQ�ׇ���^r��L�gU{
R>m���W1`���š�E�.�1'��#-i��sO��oءD�p���_�*_�!�vm�t��k~�Y������{�x���T:;�c���a����c[w�TM8h��r����yY��x�-���G7��G	��53���?�Me�A�j������H��Z8ۣ M�iC�h�ϏƯ���?铏����zX�Q��\�|��*k���8/SS�`zb?c:�}'t!�(�d����Sؙ:�\Z5�-���ۏ4�"W�����5E2���w˳�o���T�u�NQA�P�m@[��Ī�@�yS���t�7�%<>�F�v����[��KZ�[Su�����d����=Ee"^�l�m���c�3X��z����{�:0���BW. �x��$Z
c�#�c\��Υk����Ѩ/�_~�m����_M�/}�߷#wwٕ����$	��+4��D㧪��#�}d��	?l-$�Ukݛ���T����z,��1�ͫsb��N¼�pBgjsT0���-8�1/�\�xǏ���yF�:}V��yIY��´[}�ofOH%�Z��-_�?k��s���À���@쳐��X���L�i�̞#��;�t�!D��[|]��|�)��/�|��/�#s�ķ(0v��ܼ�I�k� ��s�B��8p���q�J�g�븱�H7yo�{���m�{�N�d�����)w�&�<l����3G��q�K��#]'����/���F�#H�S�	|���y;�ퟶ���|f���*ʆ/U��(��H#��Ȣ5@�����նc�������*������&�y@^���Y#	�8|�uьGan2�}��ԍ�z�a%Ѹ4Z�N٭:е��K�}
t>��ٝ���Ǌ�ё-uK ��MQ��}�㴌�}�����=�Uy������܆�[ڵs��ҷ6�"&n?�����J]{w�;�U�|#�Ϡ�?�$�3��FH�b6E=�Z��y���*��5Y`�fD[�CNS5�!�	�ʴ����j�M� �*��$����k��d��� C"�B7wT�6�}=����G�&ո���T���ei� �߻. ����y6�������^E�\��g������]��-��h,�d!	��;�[a���P��ӠV=	2@9�e:(��֞�ԥ���F<lG��<hK�&���tϛ����W]��G$��J���a��z��ETF�|����ҳW�D���r���~���nL�v���r� ���ڣ�<���2�k�m}�Ik�`������z�}/ _��}�5���7�%o���d]�i���E8�&\�d?F�����}0QR������������hXF�1)3��=mo�G{�����}��-,i0���)�P��A��v����}y(Y�
S"���o4d��>���	��T.kpa臢-�
��h���z��i�-��7��ڗ"���|K�7!�ӳ���a�ΧP�j�{�D��7�a	��C�c�bB0DC�������5���Xl=��������p�����n^��>�]�(�U`��l����,X3�����1HM�O��#($>�����$�l�d'��d���^�/��R׬�oGsm`5 k����wmԻ������ϟ_�Ar� _�6-��ύ���&���{����?����>鑏UqJ˒rϽ㒩���nΏ�Go��yv�-��
��|MOϴڔ�N��X�����/l�	}g~s�pe�������- ��K�B��/���Yx�=�Ƃ��z6�ȹD��С�;ۛ9=O��"�+k�c�PSn7-j]陸�S�����(����և��Ҟ�^����w�����tǀ����m��S?w���o�,�^��/���鄲K�m�� )4��1�PQ����EJ�T$%�E%�:����cH	E�N��nZJ@Z@bH�a I���_�����Z,�;�8g�}���2�Bû�b������3+�@v�:J2�Ƭ�0��V A��O�/NXch�N�˻�����m��؛�{<��P)���������
W��O�4Rz'�����Ĳ�*|?aEN,Y�c�r\j=���a#�6���mH�1\��~|&���|�|�LUi�e��PZ�&;�/�~�'#�+2C�}��J%��k�JSA��'[kU����E˥O=�K~�H��nn�ں�7�*3�{k��N�b�[T;�F|&d�ǹJ��_7���ȏ({�X��"X���e�>��m�K�U�J�o��F� [���Q���,�Q��g����s~W�!���>�E.,����S�L$�C� �N�VuQ��6�E���$��W���.J�9���:��	%���N�A�|ؑ�*�٬t~�[�u y�Z�����1�I���Ҕ��')�gy���}CTc����t�	;ѷ�@2:b��er["�2fF}d�8O�
D�	*0艿�s�lR�������&�*�͓ͱ'�*��W(�} �.<�^T[#��1�+�ĩk��)�K#����3l��m��-���]*I�rk��wՍ|>5��5��[����xaTNsu4[r�{~���u��NQ��91�%���Ν̷sm��?N
AI0:aږhV	g-��R�,��G�Z��:�I�D��s�s]����g��O�|Ƴe�9P��(.̥ɽy۠��.I���j,2%��5�;qxLs���*�Fk�rZ���3�2�%t3�h���^��	�֜�D��Y6|�������+�I�|֘v֠��2���^����Zʟ,Q����!�GN
9T��ms�fZ�Zw�=�1��e�YZ%�4M}7jH��~.ϲjL��"D\�Ӑ��ᷚ�b�+��	,اDÄq �idR�޽�rW-d�3�v�������WKSJr,B�d"�??*� ��w��2D�	����bjo��zCY��]��$�C�˓�����OQB-��>;eP�<��%>���]��-#���#��=Z׬F��Ȝ�s�3�3
zS�|A����&� �ٛŅP)���48(	`�cqM���wI�	�1�K��4_�ǜu�m��������v�P��Ѽ��g�n0&�f/������'�1�=7�����̈́�+3�4��	�i%�@y�6����]ňy�m��5�Pj�v�gy�
5�7r����V�G�O����\�쓝m�8����a��nac8\�	��AEw^��'�P9����A4��(�Z.L�T�/�[H�ɖ]Fڲ�D��~�a�����ߦ���!�3���d�`6"�4�X�����j�N��A���9<rr�B�N�Vb��Id!�c9�\<����B�N4P�� �:����w�!�A��U03�G��4
�(&��!�0�9 ����˼�cI&�)pU��\�喾�"ԋ��Ù��������/��X#���O��\������ϲ4wl[t�����Z�8�:����򊍝��d��jźl[�{a:o�Yɓ����/T���[�ᒭ���PV�~WZ�5{:g�핒V<�l��y؎���q��$Yx91��#�����봡36��q�z��a)��P�b��qP7E�O�1��|���ڸ���"�M��zr�J��O0��UV�&	گ����AO���)ٮI:��g9�?��qX;2�| w^oTE���6u�M�\P�f�FjO���N�&^��M|٨ �gs�0��î@�	_���g�^�ݮ�b]��6߷�����̻��Vp\GȘ�Ud������������$�j*A����mϗq\�m:rb��@7���.�ԟ��y��܆�1��Óղ�Z�L�z2�2i#����p��M���J�Y �.�`�OQ�.YjR;�xч�bL���M3ʡ"�n~B�2��R��)��V(�9�:p\m�A�8Ig��l��Đo~��f���T��j^�����*߂��Jl��٪w|×~�r=^4���1��Jj�\%�*`�/Iq�@��o�J������X���>�ri=��Di2���Lݹ�O;8J2��a7��̌鎽F��}�Z�ן����z�����˪��6��!yQW�ѡ^��ά�nK���2�$c�����M5D����7I}��lm��ق4���$s*0L(��z�>�j�C�����uגH�`�#KWZ�R��ړ��,�,f���_�͑�r����wv�a����$Hmuw2���A&O`�gcf}!��AÔ���T��~�X��Z& ��qn^�x����Rk�&\5Ae����!r�`⺂?�i�7��P�$���橲��µ�y�0Ws.N����/̷�O�h���8�%>�o��ç��)dq:K�&|ឺ�n7�ioI���o�E���8�?�P|\~���77|���isvP���Td��l�6<���jX�\!�S�+"�U@pJC��Ug��[�ٓ����۩h�zVY,�Sd&$e�e~��_?N��ۤ����V�g�W���d�>�(8���8��ˤ	�3�N4d&*��p �N��w/��0��[��$�, �k>Zb)��;-oN׎p:��ZvNP�"RwV+����8��q�0Ԛk�K��j�뻣�Q?���e�I�=��oө��0�\$M,�<C��Cp3d�?��t�"�8�a�O����%{��G
�M�[�Q��l����iمX�Y����^VLI)���n��a��x�IL�,�	���km>��>�o]�m�����֞���;����SX$���#�6Ȁ��^���Y�&9G��e%%u����;?	�wmdH<��V�Ot4j�b�
��K�b8I�J0��l��@D�w;�8��ET[�/R"��r�9sr�.�+�7C�uO�FŤ$�6�r+W���M,1��'1�®�UT����#/��/4]���'[��f|������ĜJ5�;�y�W�ae�; p������t{{i��B:��l֖W���*+�#�;��O(:xy�.�W ��2��u����g<��և�f.�6J�-���&����zT���"���ʬ�4�-y�؝U��(x)ى�%����o�=ϟ�.��n�(	�MQ꺶��hTܞj��_��b)�z�|"�ɲ�Ѡl�t�v��|ͧ>ؖ��xp����wLJD۔S`��M��Pf2jTy�>ZI5�5��d<[H�w��3�q�͏P$�Rqm?ܮ"��;�}0���> ���h��z�Bb���/.�����|�3O�3��1�k%H�f�n4��}���I3,v��D�!����DcRև���EI����<U����cˠ	}����QbQ�裍�$4(��8@�>ӣQ�fM�.�#`����a��w-pJ��k�c��A����"]Z_��#Ϫ_��d^[��q�!��r��RyA5�̬�����.!`f�tW����n�Z�� ��݁�N�������?�ղ�,u�MKʼR�m�hQ�՞g����@�����l����͟vs���j�v��_*����v�j��\��f���Z}�a�p�n�S�������x/�l310U������9�J0o�i�[�����c���^.���{��N9���>/rx#�VKP�;A(��u�g������7�P�d�O ���+�`��4��2�� xv��-�؞�Ư�i�x;��m���{ŠYUvi�>�=x�2.g��6�n�n�����6",T���a�����(:�F�q�I:�)ie�d'�����6'��.��u,f�~�<������.�v�������оq��}��Ӫ��0���~S$p�C˥˓܆ER<Zm��2�3�� 'V��W� _��1����f���k,Fv3�o�������a�/j�>���Mx����=�x���HҔK<�p��ݰ����~�����*[�v��|?>��[��U���#w�[p%IBvߕ�t󼺮5=�a�9w�o�L�[ވ�i�\�V]�9��*?7�#���8[�z��7`p�m�x�r �s|[��؇�E�i�D˷2�D@k	l$>����EY�SQ�����)��|I y���f��|�>`,��|wW�0U��׈� $[ˣI����wH֩�vw՞��3�E���^��B���#�;-n'_�Z�KD$�����{����u�u1���r�Yp$)B��˼"D�W�t
+�j�$��'�a�����`����s�$�0��!�P`w�YF�,`��9���U�?��M�p����zT"H\��g���f���\��O���N�2����T6Ӡ�g>���(�G�$|)&$���]��:��8/p���%�W^��b����菟bCwd��L~b�p�q��?e��T�C�e����_x&�"j3q��._��x@��:��)\���f�+��#�BZ�F�g�� ݏ�?�c��44�ug�aNL��=Ӌ�}��r����/h�T�VWV���t�V8�A�n ���X8���k�$�&O�<s1������w�v��F���7�A>��6�]�d��$���)JϬ&���雾��#��jJ�ȑ����� J�w1(� Ȃҹ�r��[JtJ*�ޓ�c��Tа`H���zr�bG������[f��c:�U����%�����4��S�nՌ>�X���y\=��$����Fz+��oo1Mr���0=W�m��)��x�k�&�����H�*�GL(!��EI������6ma�ک|�y�}��,�I��mZ	�Q�,�x�5��e�l�~���0�4c�K}�RB�_Zm}��}�`O�y�rK���%�b�\F=o�L�Z�F��qaޢA���B��()�TƌZٱi2M2qj,��F�
��'f�'����eƼ�S*������� �On/m�w����X��
�*����o�oLj��?��r�H �<�ƒ��>v��,��:h�)M��D��KCb�vM��o+�,I�����D�o%�<�D)�l��2���z�œ��w�I2��ZO��&���l�U��#m��_�H��"){���?�[9L�<��㻎��_����Wz��[�%"߷2 �;���Q�un�$��~�-��Y"�=�� ��r����~}�"�q���V��|��.���>'���ͽ� ����ڛ1��y�#:Cߋ-7YqW�艁M:!w�#�I:�O�Q��s�tޅ�*��Ґ5_�ww�0�D�.rԓb�{�����!s�
ǧ�'m
iz�;`u�)=l��񧶧,�/���UOѼ
�a~����a��1������Y�����C3�(E�Wƙ�r�T����N�˜I��ҟ�H�`ULj���D������GM�z���El�a��F2��Q��6��|��e�Z��N̹0�{f����f�w�O� ��M��s`�<���>�~ Lר�X������w������r�<�Pe�3l7�Ӻ������F��̗�J�r��v�K�[_���m3EZt�%�6Ƹ�Ckw�&�k�����nWL��:.(����,�[�|��lVakQ�]`����`�
O���H	nt��X�C�b15QFȠ$4�p��iK�CJ����Ȓ�������Q�F���W;�*S�Z\�hs��T���LYo��lּ�t��Q�𖍂4Ý���ґͧ��S���r���7V1)R�����{O�8nثv��D�n`�_�)ܳ׃`�l=4.�#Z*�3����s����0F��ܓ=�0�؝����/�v&�}�K)3;�Bq��Ӡ<�+ ��h����;J��$b���˓���[M�N�xtg&s<����j���H�����P��E�ͷW[(	';Y09hcj����@�IP�l�&�g���o�5T�#~�a��崙2o��T���3�޳?�����9A���Y����+f�z�W�5��Rn^?5�ᥚ։��_4��Fj��N�Vڋ{u�����R�H2��n�O\��6EF� ��Tiz>w����11����S��eM˓�-��6��x��ּ�fan��ǀn���#���11�Fa�b�4�����"<\=z'��&�~����a��/,`�>�A�)7L�ڇ�6���b����ɏC�J�͆��4��*u�bӋ�����wQj�GYwa�	$?V�a T1���Y :�r�U�O�0UZ�62 �S3�(���JV��!�d� L@y=���` �%��Ȧ�^e�oL5���UK%b�6Yq�q��\K��֭L{�ԍ�Ls�R�)��W�T��}��˕
�jl�h�m�������ݵ����f�d&� v9���WS�	��|������*��@��?n�{�*���T�Sk�W����4�isT��h�+�0�l���2.`l��H�t��z�5�|�|LBg.�lMs���V�\�j�	���%>c`�
f"/��9W���p�g�� �A�6<���aD̦P�A��u�_�&3�A
�$�F?|�H�NnGn�6�� �7���<�6��:5༠0>��_	�����'�B��C%� hB��5~�r�؛����%�!��eW�_�� b}}cסuFyr�c��,�*]F��m�La��x�����:�;��!�ڗ���p$.�zI�^��a�L̤>KM��������6#�U�K�V����[o��T��rU�EXE�ߑ�Ag=U��<'��z��]�Zm�]�H�>�IN:����t��%�� �p�<4��;Tu9��1�`TzmJ���6��i`��������7���I���;ꉏ���Y/uDCa5F�<�UK�G%��� MZm|�����q�w��ٴ˸�����n��$��3�'' С���!���+��U��<r�T���x��js���j0��<	��0�0�k"�� c�F}�vǉ�倌���-2�����~��w�S���f�Ϋ/�]�������4�\��ff����U+lGc�*�?a�i�k&q���s�9)����4���M�Ta�0� �f�2��B�[��o=1d���jR5dlj���\9���)l@��Ҩ�6$���Z�v�\��v�̀"����Īt�NB�͒�,�vz�>�LоEf��{h�!�&\r��4�|��a�@�� W��BWM�e���e�'�ڄ����c���ϧ����W�١�z]�@/�H��>���ݔ�e��#Ű
,�"�<������w�I�(@<i�#�횐��R�k�m4^�~˫a���w��c�׽s���p����B��e��%�t֟2\�a1y���T��ݩ�ds�M5x��*��G�=��OW���~�HO�S�~���p�z�\��a�Y�����G�Mߠ�0�07��p��E?b���¥9y)�?�E�HɅ�ȁ�����]p�/�o���s��^��c���y%ܲ�r�3�fAQ�|��?Z��R�9��A&�ˮ�i��xn.X��幢Y��A	x��;8V�#��l�3�z �i�&�e�Xr��_y~ф���U"5t����4S��=C��/2:�l�{d:���؞�?4�?ϯ�ez��Q����bcZ�<���T��pS	�hll!�WAr&�c�	��;�_���1�i6S��J{��w|}`��oqD
R�Y�Eq��(e��TR��d_��X憗���#�����6�|^��O���ڞ��		1���������=�����SI<������x!���%e��Oa崯��_1��"�`����zv2�����?����	�zJD>.��2ZM�O��vRHCƽ���"�I�c����\s������
�[�_�ҩ2�t󁍞njg�(�܏O�a��EF��O�MxP��z�}�7�q�����5?�-�R���k����o�)\�V���ly��=~�P�aQ�c���&�<uU�U��f+��l��n��v�9�`!�E�q�Ⱥ�:�8+nBN+3?b'�¿�՗]L:�=��}2��F�|,�rE�ʰ���1�e���i��L,K�<���w�FV������|R���"������/�W�L��LY�K�&�G��,H.��q� |]h�ev�,���2Tȑ�T���C��$��z��H9��Lf�[�!���<�����H͵�l���������:�����ƫ�I�K_��<G2Dr𑋛ȅ]��w�.��/�k���b��иͼ����O�d�Nry���OsT�`��A;Li�U$
�6���o�5��v �8wm�"���q�m�z�M���L��~�o��w#~����>�]�P�ć_˼�M_c=�!\����Z�#=ܞ��h��3�<�ě����f=��b�v�������^����5k��2���0�����ï�$`�� F�3�+N����.pP�E_�Fے����m��\��ao�nN����$u�?_{h���v����+U�(:��C<���E��t�3��`������K<�X|-y:N�j�-G��ɽR�DL:GLv��`�����ΰ��$\Ea�s�p���5z�N�g�������
I)w�oEgJ�"M����k�Xߍz�{)��@ĺ�y�%!��l����i1;�������kB�,j�?k.%��\F7Ń�=�g�PT\�E4��i5q�����{A"�nz �-1EO7.1Et��'L��FP.�"j���[�@^I��S�GsMr�j
;������L��n̳�����ޜ�2s�ޥ�	���a�	�gV����tե���^k�=ޜ�*Ϣ���ld�_zp�b��='*͜F���B!|�i�F���1i�m���1�k�n�c��җa5�o���LI�	�=6^����V;��o]�ٍi"��kӰF��)��Bs8�C�]u�L��9�K���)�yw-�!s`#D����rw������2L�Y����\u �=C�T��ȅΥ�K���2�?iƭ1�H�v2Nr 6���Q��?% P3U��v�+6�dF?`���&��{�ãH���u�8��A(L� �ܚGv��Z����H���?YA̧I�e5%4��s�}��,]���	΍ڈ�w2ة�ša|g#�+5��&�������LJg��8:���n���/�"1�n��*�Ŋa0�lww;��=֤�i?k�a��UK���B�FZnyŎE����E�L��Lӧ���^2E�:�H��R����t��L���"�v�EË���:(��of�YЌ�,�e.:)"��(��n�&�N����t7������n�ǖ�	=G�T1�*pʕ�]�s�jn��@��]���jG�iyu;�gq ��e����n ��T��r�C[�8�؇lb�f�6�tB��j5noY�3�+8���xcuʹ���#^����pn4��M
{w��E_8�4�? ��@ƽ�'��=��d���_����P˕���K��q�&?x�:�I�=��5k[����!�@{�إJ�S�JF��I,�����A�%�o���D����t���P����j`Q�M�Ƹ_��
� #�-@m.a�ED�{U?��Q��m��JB�L=�d9�Z(���
�+:�3e�����Y�M|�W�ޮk�*P�U;����N�Z�׶Eы ���o�HM��ͷ����Ƒ:Ԁ�\7�:=8_�̈́���	�� X�^��Q���_�m�+~��-:���is#)M������0:�J�����T�� ��mSk R�A�/�\�_8g�v=y&��RR��5կ���D��/3'0�/�]Ӷ@���&�`$%O
��ϳ�o�f�
���[R�	��h@B�wɃ{�,�������oH�?�*:T��y9d��糇/�?<7����>�^؉���ZfGg_�t�W����_��!�����Wr'���l�������y�	����!1��:��,e�ю�~w3EHw2�p�ձk�m����'_"�]�� Q�� a&�(@S!���url�Mn�:҆��o�|�X"��u�=g�������u��y�U��>MC���Pq�'�s��	�\���>�ք�:`��ӎ:-i���Ma��z�)���j��>%BA��F�+-��r��4M�=B:�:;ܾNfQ(���BO����DWa��%�	��7: #�8���6;h��!�����;�zF&�ϯ��ܛc8�ѼOp�Z?mh�_���l�J�CE!rU�@�Oc(���Ƕۯb�ޅ9}�뛲R�#Et�>u�&vт��=9�|�Q+��n���-�[\�����E_�Ŕ�g��Wi�d��EV���k�A2��)��L2���#;>��1v��LR��!��N;����<�WW�оi�A��{g4ל���}��K�G�J�T�j."��Cĭ0��L�~�+�E};�Q$چ�nڳۼ� �~�S��sWԛ�v~.�_�L�]}��s���fa�0ػ�U|�
���)�^�A��ea�y��E�6��|�@r�ޘ.��>��fbj}�I�{_��H�>zz�,u?,W^ڇ8���<�;d�gƅ4�6Z[�#�z�V)����]�r�R��5~�le�T�٪A�0W���Y�L��T\D�=;��gyW�̍ޮ�7��2��u�PEI��}=�)�)�`d2�dO��d�j��V��U�����OZƩmȰ��QW?���Ih�ݲ������?��x�*�Oh�,��JEӉEe�����ĕ�&�L����l7�B�|��E��Z8�1��L=�JY�e��cܭ
.a�1.�}D���h��<L�W���ə�@W�U��uyA���i�5T�aN�˃�&�����VG����*w�2b̒��we�-�GÇv�zn�j2�=/�{zWx���5��N�IB�oOf�w�٨�J��	�U���q�Hb�ԃ�!�j�o�.��V����qFv_6"
��?>b���g3~8f u�#F����g��/�=׏=�w# ���i��i��d�l��As������C?��U�:�����~����F�	]��_�\F��y&�Kx2�����3Śi��py-ə��7��Y>�y�1^	yAm��ƹy��EG���Y��Q�/By7b���Zt5��%-��Ӵ��J���[)����y�����������4�M��eJ-耫F6?z������^�v���^�{�L��vm��M���3�ӧG���ʇ��Ȥ�w9$#�*z=�̍���L���o��Fy8��s_V�V6�%��@�=l� �,a���24���������\g6D���y�������ڗ6E�h,�Ψ��&1�}7b.�iOGj��,��PZu;}*����{�<0��=x����!��7��~���Æ�5{n���o��$��ظ��d�vV;�i�M�����hx�n.�i�����5E!zt���D��� �(����"/�n������SNk���ϚvU�bԝ�v>��)B~HC�E�"}%0pYj���Q���a���^}�ٸ����}�|9^��J��׉0��>���;�������Q�n�tCbz�:�[���Wڵ6��,�g�1������i���ʸ��$���n�&�`��:<�^�[�L<O�SY��T��pp>��_�E?l<�����l�?� d�6�.!񓥀�����>H	�������j�7����ǒK�1٪�B?��*�V;}؀]`�|)<�;��3������>~/v�2�+�n�o<c��	p��QVW@��\!aa*�L~#T��4t'¹� ��u�ћnm�yol{��)�#t �dں�F��������7�����r.޷�8���E}�+r+�p���aސ���d
�o%V�[�+s�$�M��#��4��D��������M&�Ha�S`cS�>�_ 
�IK���N���>�$��}�mwQ{��u^��	<��Z��&<�os*74zq�N=��pՠo������9��7����5ɖ���ڳapحH.��|���?=�����v9J ��U�{cV�\�^�4�cC�����ݪ�}+�/���1��I���m����@���Ta�(�`6xb�q� ��)����̄z�/���=	��G��j�`³."��&~����"���J7��߀5Y����8���Xy�A˱��A����N\
xӝDn�dbXT��m�V:3Us�7$�TQ5B��x��<�o�Tb���G��a[�n`�|-����|����V��r���Yu��|�9���w�&e�g�[�0p��9�|�s��_Q4�0�T�О`�WU ��P~�&�~#�bcbm,�A���}����ٓf�a��?փ�Ε4Qp�(�Ь㇊���R�ذ�7���c�r��R�d|a+,�iÚ�����h�l#�¥@��|�@lm��\��Ll'��?"ur�;��E
'��x��X��C�鿡[��ו�ƾ
�a6���z�� Bł[[cb�h0�;�+8�<4�_���1[V#�HW�����\�awf�o;��re[����/�J�lՋB��ҵ\	w{5��E���f��4M�X�c�o�\��'iH'M��p1����@��W(Ŭ.�V�b���Q`([��/�jx�y�嗹�SC���b�=K8���f�ьN��R4
�`���U��NBρv�P�m�z;zUȶ����숏�z>T�=9���8�¼T�2���?��n�'L����Cu��<j����R�l�c����F: 0Ա�F��̍�l M�S��L�7R�Շ1S_��ex��<a����A���GBV�{�����<��ĕ6B�K��-��R��3)�ŷ�۟��,Ƀ�J`.��\#�kz��j���eN|��
έ	yS>�����Κ-�3���gh5��)�9qʛ���������ˑ'`�X�����&MbeMZ�z ���\����lh{�s��MF�*+G7�7������D@���2�g20w�Xod��)�h��b~�Ø�B�Y*�-��2Iڡu��;���Vt���Y�(��@�L�f�����ZpNr��Ç���V�Ig]�jV,��c��~��ޟH=��������U�^4PD�&��d�s�e�o/��3hX����%�ދ}x �bht7J�F��*oɅ��T?���G�K�"ҋb,�R�$j�E����Л�!��Ոi�=�M���YV�ڋ��>�s�W����h�悄��E+6xQ!��}��L�����E�kg�r�;��kE -� W�Dw=a��N��Q��c�!V���Ӓ2�|�la%MF14�0lz�Ј�6�YG���'�H����l�0XHr�m�S�Mj�!��^~��MFf�39���ظ<����g��I�("�A���s�&x�D~t�&	�O IE�������R��b|6J}��Z�V�f�۽Ql܅���/�C�m'�FP��e:et,����V�a\�-
H�rp�A`Q�m�d����(��XD�o$Od5O0U�,���k}Ƀs���sko��99���� ���y�Ǘy���[�ϭ_�zӘ�FC|���c���r��gMl�N�]Pq�RF4��o/�꙱�:
���(pg'�2�BH��x�Ɠ�4���V�n���9h�T4ʉ��w���׎k��!t/�S8�M#����}qAseR�=]�7Ɩ��H#hJ}�i�#;Rk�h�7WB���`Pu�G�J�E|[&���v���ڼ���뫑CIc2�[ZZ������%�����-�r#]�!/���X��j��,Gy��� ���+���	�o`AK|^'�:���g�ﻎՄ��J .v �\��s{�_�����6<#B��8���_�̶jt��E��].�z�Gb��s��凴T!���)�B?�n��H~ֽ�� =�p�B�b�BK��\��%�;��֯ ���Ϧ�B_����_E@mcyJ�fj?"�F1��A�A4��V-�X)�w2���Z]��J&���8�B��X&��z���4H��Sb�&>W'9��+��b
�Y/1��nzsv��ȿ)/�f��Ü��ߥ�ʛ� b	A$�RN�����ۏ��9+5��ԁzj�P��8�Y�LJǠ�)��<�J~<lK�Q6@q	]ua��v�u
����z���>oO��]�?wg����
B�I���b�©1�7�b���f~&O.}��*c(�$ާ!ĩ8i "m7T��K� ��q���Bct��R���D����dJ�p>������;���R�̕_b΅A����y?P,*�O��+��^cË�i(%�m��i�v��H]�Ѵ�"H_7��$Jй;���X�|�Q(������@��Cnk�j�s��L�9O�����3�SG�h�VV�q�E~���T�D��$�B�'��[ �T��G�GWIx�T[$Ƃ��wK�R)~����=~B�A�
��ۨ�����]MS�m̱J��[�ß������s�}aX�vt��F��>�	QS���,���u��g��[�ߝ&od���f��~�W$�L=b(6;
�R�hfQ��ג�b��VvŔ��r��
���Y+�|m��=l�B����e��w��cğ���ɨ��|��Z'�����+���P���Qj jb���+��@�Gu%���7����?�x���l�#���xzC�𣍕W�/G� �;rd8pn����c�����䋩�j�Uy��K&v��������o{�:�{�<�hq���Q,�;��\A����X۟��_M�,�J�����?sVTN��Qd��\���#�%,����db0�T̟>Z�JlH֕�X�&�Ҡ�BE�%��?��	��f��>@-�N�I
��[IFlp���kh�X�f����ۆA�����#d����8���H�T���gEy����c-D�����	w�T�"�agc�`�<�0��j��h�5���<��ˏϜ�kF�ۡe���p,�e�G����I+�yl�k�柑 �����g�����/�s�}��T#��.��GE�O��`��į��e�F��1�֌p"��Nl���7��Dx�w�j+��`��Q覐�l�X]�'�Go(�+o�<����%x�h?���<�YՠMZN�9Š�9�;ܷ8�)�WE�9\��pAu�P|�l���?z�yu��FP���n��ׁ��;XK��OZ��ip�����s��f0��:a����$���{(G��}�u|$�˿҃����{������#h�6֛`-��u�N>~�[Tv���A�t�l%�������E٨rB��ZS�������g�1p��Σ��T����訤�9A�G�N��ȎQ� �#�� �<$��}	ƴ�i�پ۽�3M+�w�"�x���l����|~~��e�:J{sG��4R�du�Հ�~��";����)e�2��Q��@�r}�>uǐ����1w����G=�u���&�<gg2W2��q{[�ß���¹���#�mV�?2��c=�3ɽ��O�
�q����b�6\���]{y�124A%8r	��**���t�S����۾���jTmnm���9}���Ӥ�Ҁ�S���T�K�!}�|[w�t 	�BL�����44��S�Ό<p|�~�
��7�ȟ�����r��HO�E��y7oq�ȳ�N��%�[4*�`ᣳ�he���Akߥg�����`�H^~���<�ʳ�/�f
h����d9����\�3AA ��ڔ P�x`p	��7�9[KNy1厓�<zsp��la��'M�od�>PQE��p��Go/}3Zug��<LOP��zBˣ.�����t؟4k��_�l�4�5
�j�fo�l�
��X�A+b����g_욺�|��ۓҨ�������!�8x�3C+���]�ჽ��U�'L���!���v�ѥL#�_hn �-����xk	.���ʒ�ң�?�w�]^�j�k��.��8����n���i\�_U�P/s��GQN�d@��A�ord��bx ���7a�����+�k�{$��V������K��?�*��2��`W�w*�F�'��Ծ��Y�ϰ,�A}��Y�*���ᾭ��`#��2��eT4s?��(�)K�&#�ͯoo�-5R{m�髥�8���7�8n�F�$�Z�ܪ�T��K	mu�T����]���mk�#��\[6��?#$�ّ���JTm�#�ԄQ�����R�P�:fhG��wR+�|E��a��.�;�:�>�\�����X{	`��b���y��-��d"\H��O0�M@E����!^��z�{s�4�)���ֈ���SNX�u����,:��5�-�� �r���)��6�������J_�1P�}��4�*�zb�@��y>�@1g0^�͛��xh`F\��#���Ja��U�����,Ln�eaiкO���x#qA���ٿP�Ck�8<��5�3��|���j������C���Qn�5��K��u�W���z��~$��fT�.x4~�ߘIF
#� �:�GexF����T�����:_�=�,z�"!oA��U��#�i+?H��X�B���������UA��1	zR�!���.����z�o�z��K]]�bB6�#4o��w��B�W�<���x�'E4Ъ4��y|�1�y�����k����1�b����t���L��)jN��s�|`�}%`�������/�u��X�2��P��TBe�JM�L��'��}�x��TRK��%GY�[�ě�o�09}6c��u�NשG�X̻3�Ul��eV���T���!�����\>�c��d�hZc�6��O���CZF`9T,ɉ>p�S��7G�J�}����R.�j�Y�$��糰U�ކ����L�XY.��0�� Ы�l4����������|G�'���5��ۗ}e��c� 
��;�m�d�n-��` �mK���p?�:����nj�d��5<́��yOv���������-�jn�� �*������;����/WQ��RU��ޫ��H�A�Nh�G�T zE�4i��"B@z/	E��w���~���y2�̞��^{�I(��O=���yixУvk���QXP�ԸWf�?}Lz�b�s�ս�㞾��ob& `�_<��B�j<x���	"{�9�ny�à�s�~JrjM�Ζ���V���+7���\&�/q���D9������mؘ]%$��r~#T?tM@������jN;π��׾��{.?�P�(��դ�#��[W��gd1����㒼0���	���)��T<}_4#���!WB��X��LC�&����O��N*tCh�n7Z:[]\#�y�O��p}�����Re85N�B��ܗ͵�e�,��6�4�I�;���?��.VKq�ݻ��$T,gdD5b�od#?�r��w���V}o�A�Kg%�6����n��O;��3��L���G�H}��~�4�����̉����`o���&h�+"lw<W�߬T�U�#�$���t�� �m5��n�&��rLk(_'�n��{�#>B�'��~CM�����t�5�gX4�OuUҋ�<��y�ڱ:8z�ߜ�4��j�Է�w2[JR����D����<��
���c`�Ľ��ϣ���t�|��	��5�4���BP��w4���{v�'9����s����5Y,��Ui�H��(���v4��p��FC�Ê<����ľ����ܦ����'*�]8?�sEf�x	�_Qmm�Ѕ)�x�f�)H�oz	���9Y�(*�R&* &_����c-�]}��L�x=�|s�x�%͒�I�eIK�=bP�����o�kz���kDWsZY�����"Z�p|׃)�^`�*�a��x�!P0z�n�;�����te�ZW9	����Ҹ)��!���(���ë���u	"�<�Gv�+��si�-�V7���t����cE�w�I�@^c�!�D���Yrb��zkZ��o�W/d�}��k=%��U��dpV��T�M�L��(��pd
���:�� �$��� �b�@'u��__/�L[���� ��D��2���`�����?���)��~0rm��P8d�)h^�Ͷ$�ڎ�o���&2�ٵ<2N�i���,���AF+G�a��gU����S�-m���x���2|\�j;�y�G~a�r�,�G��$<c_���cCC�*���	F��,����e����(;|f������z�h[03��K����k����Fo��L4��2�Wv�Z�����6?�/벷�AE��u���RA�o(m��S��\�%{sT�p%�mH�$����{��X^:[�(r4r�������7S(=�$G�@����������ƥM,�<rbxIG~rv�#=k��+�"���D|2y��X��t��%��4�,b�csEFs���jC������3Q`���Y�Ӊ��3�	������hl$���I��\�PVШ���!�/W��`���O���ݣ����O�7v�t:���D\�dq���t�$�~F����vF�9�c�~��?��l�h�Ŝ�O�t�sR��>�9��as�5,���%zbP|�i���Y1���]�viL��zmV��\�Έ����]ۺ^�Y�@u�lv�q?*8!u��s>�9X	�^+<X(y��I���<0Wr�Q(��Ö�mV�����M,b��c��(�}����ũ�%�k�lv���%!�D?U�4΅Y���r�����5�$������7���U�?g�X�df����;�m;�|}�dz.JA/����B ���9�f��M�O\FJ�w]��L{~+��U�[�
8��h��
c3���\�ޕٱt,T�f��Q{�+�_��DMρ�%����ܬ�x3�]��?�=pV]XX�zT���TF]��$Rj�G���1��[�ͤ)��`�{s�c��_��3�k�����RX����w���]��[`����h"H`�+�����V�u'��բ���A{C���P�!%��9o{Ô�f���>~�5�}"x%�����*�����6s��|�>���^ۤ`!^{e��q����X�������w���F
��]��=���s ǜgD�]p�\�{JfN�`�ڣ�v�B��SVȈ�5��{�{'n{�7e�0^a������ �9>���AG�8�������Щ��:��F�Zp�j��Z�ǵƒ��K�g8��U�Eڰ��P�Z��KF^y�|�w璜�v��nE����))0��L*F)f�
\D���ϭ7ז�������?]Y�jG��]OuY}LL軣7�Q���qM[��|�*���1#y�s�l��of�������/��xs��t�6�}?�4@��]��tDsA�Z����e��I��`W�e${�n׬��pG��5�шKz�?}W�]��9�~u 
}���,:�X&g�JhD�����j�iQT�u������4���V�&e�פ�<�|��=��xV���x��n{��k�z�<:Y
��>��vq"����ߊn9��=�x�xg,�bʍ�ԾKs��@	+�Eb!Z�H �|�� �Sa&j�.�)6��k����s�v�QF�I����c[2Qm���%���.�x���L�Z�������`�Wy�N_sY���K>:�;����;{8o�c�gB�V�`���Mn�/��>�.d����	��i�춇w��0I�(�8�'zi�(LDS�\�t���n��
q�L�x�f[V�r oMoD-f���$�N��wCE��_�=���c���גA��~��"C{�ֶ��x��n�;
�8ݖ�e��е��X��i��P䝋`�gqz�ۗ@ܱy3���+����b���G\	E?j3M��/��ؒ�X�N���M��$H&sj�)��CI������:��J�E�U;KW?}��"N�K<��#DM�9t\�Q6k���yEy�Pѕ����?r�M��t��Di
v\��ʘ:R<vM�Ρ������>>u7����o�%������
3L��������~�����1��m&13��w�s��mI!I�nMD9�a�q'q���Ω�ß�fឤ�p���u�'lTJ�ns� ��/w�9��*�%;��G�NUR��J僎���\�86���jSK�N"�S����Sow��N��2'<����mL g�z����`9�R�]6�w_���������uFF��8�M����������bɴ��i'C����D�ݺ�T��؃oa:��oVE�|
�jiy�����Xj���]� L�6n�&e��5��?J���W��2�\Jn��	�3@c�6M��X<�hz������T�;�R����Y�P�G��j��z^T�⃟�+Wr=������P���Fr�Ȧ�� �
n�st�<?�?v��"��p���R�F��#eV��	mDW�˳Fl5&�
�t��wY����63Ұ�4l�{Q���:,����,�ꘈ[h��O`9p^i���詷�w�Q���;/kW9����?�o��o�-?���Z��YK9
���w�4�%k���ޅ�b쏵-����8�T�}���ؠs*Ǟ��pk`�`c�Bi�Z�(�Q�M�k��|��ڽ�!�ֽhU�� ��G���e�u��F[��sO�����)�O(a?5��"ʑ3,��J�+�����Y�(݉�e��q���3�y����3�Md�	+6��������$`ˋ�����
��_��X�>�T�,�/3��+0���/ �5j�QKK��77 ^�ċ!����d�ib��������>\U�U����z��~~L�q!�$���bX����ȫb|�W.Y��K��l�V�F� � ,��U#h�iN�+�b�I~�8LւX�=��s1�c�Ε�x3P�8��.�����p�ی������ �5�;M��
�*2��LWW��d�9?Ǯ���>hY��2�E�N�H�q~d����y�y�k�K�gE����#b� M��6Y�	��HhsXJ^bwI-*�y�T����G79�� �{� 5y�в�#�-�d�0��c��ݳq��5Z���>I��E�I��Rp1�d�k��?�[�]D9'��$��=P4�E��K�۷�w�����r12�w{��E���r���J&cQ+#'hnȤu�(�[�jS���哓��Io�2,�%��SfK�'�86نĄ�= �9J�a"���>_;�v!��P���K
��O�|a�;��9��l���T����|�%�L8�C��ޤ��1<�"DgسD�T'�$�W��B��z���1���F�����ҎPx�4��/����'!���-r��-�����&���	� 4_<{�*0����ݥ�
�Z��(�|Vj �t�����Z,s�l�1��¡
e�Z���gM<��ߟ��$>b� �8(*�˓_�mHUq�ځ�J2����5��u���T��ng1�Ax�j33����fف�~R�l�x�<70!��z'�5U�ͧY!�T(�T-o���I:i��Q.��g%j/^=��
��K�)��r-6l�B���GU�ϸ85������*���:)Ѹ1`w�6$�Ѻ~���x�Z[?��ʈ���y �����k��s��UG�~��f����F0�a��s7��*8�#\I4��[V'�W�B���BP��qFK���46ӳ��ӗI��v9@�F��Q�K�o��W���&O���B
v6 <�eQ�����~��0_�7�d~�9���]�Ĵ�U�Ѧ��w��}K�������k��2)�^��.!Nz2*	���*&�rl��!�)؟`��B{�#�}PG�8�ݔ�z��e���CRc���}q=U�}�9�)�����6�	��w-�:OV���������l|s�	�|)#t</���k'a�K��f�-DeS44
ٙz�3�L{�<�xn�y�-������"�����h'���������t܄�.j�Jh��[o`~Y9n�T*!+�Gd��8B83`l#�`���l�{���a��o؅'u�5�w�>��Z������5�;M�5*Ю�=�L�3Ԃ�������t���+�=���?�F����%�Wn�8QϢ{���s|�A5�FnI;Iҗ!�����Vn�49F/����X�b*Z��|K����~�N�@S��[靟�~���i_؂�G䧖��`�� �Bu������~�^y�mfT㗈3Q�� �����s��>���AH�a�ǫ-�K�i�n����5�Y�tIzq�0���mt/_�S�T���7�W��I�� �X�t���<(1IDԝ�dZn�߅$5�V��S�^m�!V}�3��o4M��~\��k�p�˿-]�����=�r�$��" ���_JW
p�)G@�3�$�AA�ڂ9���BCbO�t����T.t�{�Z��"����z�P�Icz�Px�ai�}8���^A�ᅺ��N���q�E@����z�х
�@�WooYe�$��$�xD�nߴ\���FZ�d���KVYn��-b$���=HS�iS�n����,����|��	��hKi��d���fX��9�ͥ���x�^%��:��!E�M~��������sx] 2pX~3}��-'8L᝻$U�RuUOuU�9�i�S�ɾ;W��Ia���c�U}˝o�#��]#g��N�W�Xg�ˊhVMv��$R-�]	9w�������] P�^�ɖ��v�9�*͛%���x�砻|d5�k	��v�����ߥ(��3�<:��r�|��_yyS��/�KA"�O����6������f9�fR��n�$ͯb1j\��@��g"sQ�Y�j:Z�Z
a�Ӡ[r����hf�8�6�"�a��|7��K��c�o{�d���s���g۶|N�	�^$PJ�%k-l�NB�� �a�EY÷�1���+a����+ulGɻ���n�}H:���� �I�A�0���W�-4� w�T(qx	T�~cI�Z��j��UCvu|�1�p��셝	Jdꫲ%�4Y��l�}���U��F٤-��|k����ę|�k^9��Qվ��=�g����caX���];��L�:�0��07
<n!�W�Rr{��Oԛ�
�9����J*���N����
��hD��y
��a���qӠ�B�h���N�����؀�����.�"�f����(�~%�FN-*�����������oMB��UH�q/]�?U�n^S���CU:ۇ�V�;��=B�dUXEf��T�"EZg'�nz�N/1��p��0�U�E\�tS��x�����%j����=�W�ɡ���]��)��iܭ�f��d2��8i�Os��D�E�a6�}���u�U2��BS����n&N�6���[�=o��*v�,?:ό��;s�[�2`�F4��l����A��h�t���9r�bS�p�&^s��U�2/��ԌЄ���_R&G�����K����S�xʉ���>�Z�)P]'h����kP��� R�/�BNY�N�W���'-K�M�hb�����h�/i���+�Ԍ?x�� �2�2)��"Z��>���a:���Vj�����&��oSh;W[.���Δ�v�y���.r�͓�sZ��޷W�»�{^�p	r~r�:7�M���.鏱����J2G���Qg<�k��X�fNXv�KJ� N&��y>|5��
t,d� �<s��"��:�Srx�<��t}>5YBB�4X�5Ys����]��C)X���B�;. ���,mǕf�l���"� ��\`&z_]m~�I�P�s�	�f\�P�t��z
����E���xnWH���d��#�����e��*1!o���u+�}"��U/cB�ɣ,2�B��>���5�a��}39�����X�f���ܨ�(��w�OI��3�����Gd�Y���~��!�F���*����BĽ�_ߝ�8��3������G��O�?�F��f��y�6$ ��qvh
�f.��e�B��tab�܂f�UP���ha�g��!q�/���Rw[�@e�w����a}z��q��I7��r���)�DG��f��f��VAWC9>����\�	�죇��g�1᳁�y�[>����:;�E\��u�V���EX�D*�i�"7F�w�y���#��Lvh�銽��NI�z��)ߝxu�]��F��U&U�mcZ/����J�_R"�F��Di��u�*��������˂���9:{�u�~��R��t����=���Ȫ0�{���",�!k��'�܁��4:6[�7�6S���2��'hm��3�^������ޱ�Go�Aċ/ƞ�c��9�`9�*a�y�L��6F?� <�[£�N^�LW`�[l��i��V���\������}S�����%O2%�J��Da��}��OX��^�a",�Gr�Y����.�%�	ǈ#݀�q�?��lNZtYlRH(�oa��Q��&��D)Q4�Ќjggpj=ŋ��w�T���ٙ�Ĕ�}������\�e�v�g���L����"غ�HFV-o�P�e�8=,��}������8���ҋ�ޛ8%t�ړ��.�~�����v������=�_�)����^��f2F��/O	��ge��V����t�%�v�F�I�8��EJ翪eD�$E��Qε������F�^�!�W��bXH�n�?ɹۛ|PФ|�N3S'�1�:^mB�]��D������Kw��+�_R����U9�f�(��џ-�u��K��BC��i�'���������e���59+M?�LxS�
I��%�ُ	����H��ݵ���	��R�K�i�@~r4�Ƈ �ۊu�����^V���'ޢe�>��������P|�B>ȟ8��x���y��ni�{�,��	Y�:ʢ���H�kFr�VG�Z�\}�4ת52�$������9��E�MM;Q���#��>Q:��\4��Cq4��ɗ|���\��,�m�3@�g���La����7�{��h�l��Ğ��M�(l��/�(/Z:-�k� S�MFLsz�_��"n�+�~��iA�H��^�!
X
V��h�%KI)�(����{m��3䝧Z����C���M뜄���(2P_H�������$�x�L������1��!�5;9��&
吨o<X�:J��Z��� ���:"_��Tvv�9g	��I��>�ٝ/���B��g^s{�k�^J���	�c�鞛�q�d10��L��
�>)?)}y�4���l7���97���4���O��"��jt���p9J$�yS�YW�,Z��E)�v��ZD�����4>���s8i&Gj�UЂQ��i���7��v<��D��
9��YU�U¹8��C;�V���.�l��x��9I�N�5���x��L���a�K[	�g���ӵ-[�\�؉^e&r�7�:��dj�>�$�k�9��u��P[�*���L�w��	�w6��}�֟. ro*���F�;R����틆�~�tf�)��Is�����Xs�9���� j�mZb���}��}��́F�%��E�7�AZ^��_�w�@�P~Yc�c��"��x-�W�L��⟃���P\Oy��QcN�1_�1Ꭻ�!_ɐ�e\Pȍ���Y�������J�L�eB>d��З�Y��<'���Q��R�E���RCx�ʘ^��φ;���믦6�g��4Nպw������e���೸��|pP�8M^���4B����?�/P�A|�Z����4{_�JᎽ��U9�:(���Zv���(�o�<(���h"p; ��	pԯ����Q�B��7�gLx/�l�Q�Q�9_+A�?��}C�8��/��XwśR�"��� ���a��Ϛc.J9�>/����Q(�"���!&}wAv����;$��m��YA���1;�����6��p�='e��	D�.S�x2�e�1�滣r�sLô7��[2�e��~ma0��m':# ��t7�r���%�n|�g%�ӛ�+RͼAР@��UϚ�ǌ���T_K����ltL��|�,��<���<�#���/TS�1R�Wf����k�E�\�P=�9٨�;K��^��hp���������a'EЈ�A��;0���ef�M�}��b����$�i��u����yf7{dܿa���R�_MIZQ���^�k�Q��,@����oXk���۝Z>��W�y|�qz'-����QE@�`8@�"w��X��D*h�s1�^}�aL�'�#�<m�o���&�-�F�.�&e��8^�B�T=g�;8��F�=ޔA;�S��,B$)�u�}�%�g'WN���M��ٗt�ܡ���D�M֟���V��j�׵�&owyb�V\&Xu�T������iGe����cɅPXO���f�^�	��M�YZms���2�-R^Ұ@��F't?��X������mۑ}ό-`$)@I����ԝS���M��7��ޛ$�(fm� ��u���=�y�8�} #]@r�%���`x�`%PeNV/�'O ���sOƴn-y��\�I�r��P�i~�aW̲Ȉ���L*W�ќ}�ʬ������FԸ�C�Kɮ��8'kMc�3�/��XWg"�j�r^��5c��q�gX��qU-7� ���"T��,|����*�^��Sy@���k�'�u<q����)l�>�q1�&Q�������b=����>��I�,b8����|�fx�\��ɽ�gO�<�
C�N���ǽ^G1���צ�OP;Hl�A�ǥv����ƻ�h5�h��E�2���
ϸ�Ҟ��f�v���) �x�ʹ]��wx�P)7��:r�5֋�����j��pz2�2�\RN��v4n�%{��>��>n��O�j�͜W�5ڽ�Y�n�M��������	%��h�T٬���E�sŮ�p�"�r0�[�u�7kɻ�r>���wCT+Ww�;S�[��D�zX���	;�����s8浹ö�ɠ_�˳������O	��w��.�~��s��2�9���H����x!z�)6�l4HY�I�#�7�PK   J�XF��-$  ($  /   images/d88a5b0e-66b3-4edb-b452-47f46dd40326.png($�ۉPNG

   IHDR   d   o   %e�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  #�IDATx��}y���/+�ξ�o��[-��I�,�as�k�k{b����Ĭ���X�ځ=�����zc<�'^cds�!�!	��VK�-�}TwuY���<��ZjI�T���̪���z�|��}��p�����>on���,?�aW���Gy瓜{��گg��ש}�w����7@�tvT��2 ]��|j룰dO�f�>�}[)uP)�{���B����ත����0ۂ���G"�[�UEoUѡ
:#N���@l��Ӵ?�(��d6��F"t�"W�� ��b�rR���.(@޼~��`BS��i��b-'N�$�^G���L�&�m#���X�%O;��e��"�>��$<��v']g��/9��ou���	S��;/��!~ d*0I42q�C1q�b)��Jb�:%&�2�J�#=�N )q�Ɖ���]H��U�Oeo}s�����؂�8�ca$2!�>tp� ��.6l�`d��i�,��b��L���dSv%���ޭ�<�[�ʲ��߲JBj
A����c���cy��<����f\C�`MC$&�SI�B�{M�W����}�o*�Q;�й\������u.\�3��f΀V�1?����rȆM>������� �K"��f�⿧8t�R�<[:��ZjtN�H�'�P�N�0�C(�A/��M�6u`�z<'��.jF��R�4R{��8"P���F*�h��R��w�]\G7AO+���rC$�r��;�)��� �q����wl 9���iʠ����0��ފޗ�";���N߃��/C��Q�(�-y/�N=��ڊ��6$��3�f�C_K5�,E��-��Ș�5I���������9C�5���
����)ddK��@(.0����bٗ��Cli=�<�i�������М�pB�B0��;g,��`dd���+uZE��Ɇ���/�=�܃E�!�a6��+���v�F�2�B� #�����l{�3�$�1嘪�H�QT��	WR�@���b��4h�-�|~�, c�0ad0��1Z�@J�Ĥ���0���*!�?���� d�-alղfԮhE�D���C�X\�ٜ0J*���͛��s�!�N��c�Nk�o��F|�K_B�|yfh>��v���}��R�����8Z?N�������]�1����%Ʒ�ёhFk��^W�� �B��r���e�H��5h�$���z�C����L��.�1��O����l`X���9��Ha�PV�ԡ"������J�q�X�|9�|�I������S�r�J|�+_��^t,
A�4y
���0=��a�X��oB*�'a3�t��4P�����XVَ%��D�S#"):�`��I��҇�e� ���J�W��0�8�@�����V"g�W�ƞ�c�=މ��0g���
��3����2X�]�yÕ����y���_��9o�<|�k_�O<����3$�s��8�&����Aqm��݋��QX��.���o܌�<�l���0�e��Oh�ê�K�&�X$��ּ���3�"1�\��LW����A	a�z�P���0�H(���z,�h�����L���Ǯ�Q��aE�*���8�2LDt���>�0�g����P�!444�z���6�7�,,��ߎ_��gȲe����^tQ����_��ub��M�/@�|Ri����`�s-@�D�$���~	��,����#U�0\�pU�H@��[]�� ��baK����*��h�8�f,�h�p�������J��a��}}"�?84g#������O�{<����a�?~����k��/��&&&�Fz�t�k��@����������x�w;j��9�(dl��>�6 �>3����+��v�HG��E_~��H! F�Ĝ�J��n$�¶> aEP�!��v2�`��h�J���wJ�(dD�B����1�t���+�������7����G��v�څC����ڵk=PX}%�I�T���wf�TWW�pVSo�����"��/~��5�nˡm�'ȵ-@0L�=u�`&�^]��hX�d�R~(��,�s���$!�խ�
�3�S���H�-3�� j �WJ@��Q�φ�*�(�l�W%����-�:v@���p
�<��	��_�Ǟ��z6��<ۍ�����7�)��}�Y���<�0����3�<#^ß|�OP���I^��y@��yCGC��5]������dq��h��9�
ny� ���X.(��*O	=�+�5�A0lU�����4r���*ɵ�Ӷ۰���3�o���s�{̠u�i*.{�������-ro�\��c����sp�+=#@�����Ν;1<<�U�yU��8�0����v�G�0�"0\�}y�"|�i�0�??�4��'0E�x�Q��#n�0��3�;��WB�I�FĴ��[1$O[�uqUǥU�yh���%6�>�cAàW��Gn�B�����<����cŊ�<�3d*�7Ŵ���6��a�Z�9W2�@ gmf��WaUr!�I=�D:X%�De�gC�*��|=9�E฀ؒ� ��{�dDD:t�W�ለ-㇤R��+m�`���7���d�\P�.���M0���w�?�B̆f�A_444$�s�Z�䟮��gUe���w����-ע�\���� �f0� J^�q���\Ȏl�-g�*͕���+�tn1+,@��QS}o����VH���/�'Ɵ�.�.����$��,N<�'N�Άf�}2��5���[��E� �i8@����^ppw��� �m�8��D�i�t��������F��)��OM��CgUE@��߆�ߪ�[9�������v���� ��:���C"�\N���Ff0=cw�T� ����~)���<
8�������L��x����'s��dLP�5A�-�XE��.�(�NݿxyF��P�,4�j2\��u܃�s��<9]�iX�������N���K���+�_���Ӌ��-ۀ��z�=�Z�[�RHQ�́���
�D̆l`���U%�����T�׫�*��w�GǞ�Q a���M�����~ؐ��贀�t��u�U��� ��au�6���;Z�̏a���ƀ0X��'q�3���4ޚ�tx�n����I�λOvn�	�
v	GZ�wL�汫uk����销0��k���4J�e�)�Nus
��s���'?}D���p��B#H,%�az�S���T�P��fP�w;���g�!L��`wJ:=�Ćͣh�cA:y��90�+f��k��3�@�QW+�pK�:D԰dL���'Ĉ�b&b5�^�Lh����)��H���[D}��80epD�jߠ��1�p�)�dF@�wmO���Y���p�aUuC�*��jě�S!@X�ݛ�(��խ�S9=KL�p�3��������o@���$}?�OG�5��{gd 1���r����{���K��I:a�����^�ǍX-�������I$;`��Oԯ�k��A��÷'�%>ܘ�Puι��thF@N�PPE���
V[qԺ�~�H����Xe��hy���d����M�s�-7�s�O�@q���5~�B�����`*	H�MKP������n�*k]�R�J�s����V�E93G2ܤ�jؠ4�kpϜk��]/�t��K��J���������= <�u�c���~�?�����X��K4an�A\���<P@�}/��ڙeڎ)i�o=�]�������t,z�l:h6r)V�3� p_B�ĕ߹��]GQ���~�ignY,W&/!�v��k�/&b���?���%CR���Y��tv5_��n��X��n�Q0P�����w]G ��M�������"Z�/Y2���p�y��%��jQ�����XSx���%C2ʦ�Q�TQ{������N�Ԑ��آ��!����}������0^��om@b2'�bZt-��b��C�6N�Z1�c�Q�3>�Ĥk34�����t~�q箆����>v@��cM��n%0���v#��
 �R�Ib��@y�1�:=���(fR"��E���g���n�F�{fM�Z��^��Fv�"E��
���3z�=�u�[yK6K�G�!���n����l�l&7%��b�%6��k��*��"NcЮ�[�w��;���'%��|F	)���S���]˲�.��M��ڽ�q�'P'��K��dGܱer(�0=bp���awK�"%<�rab.���U�SAi�<}|#�V�`�4���>k���=��rs�n�U�t2%ŒG֑[]�wh�îH.�މ�"%��(,WF,|����y/��������@Ϙ�{�"��0��e0J���H_2���&/�l�A�,1�'tM�3q�PH�"��5>@�b�iY�f0g���$t��q
r���w��/[�Շ��(ъm�q�C߸{jk]�M�y*��52u[�t�2�����!�2�̲%$�-6˫:	׽�Y�U��v��r�<��k]C�\pF��1�h�S�H�3����Ɇ���<�I���$�rVY��V$	����<n0�#Gx��L�,�i�`9�@�}�}VcI�!ܑՕ���&��d����I�%D�i��n�9E�R�fG���c; ܑ���T}{���>?��H��w	���"�0P߰��rg��ivda���-�sj�v����r6���i�Aol��Z���*�8�a��r@��G>6E������9R��&@��A�p�?��0E�e<Ό$��p��w�Wk2 �՚�a10�`��,!��l'���g��9sr�(8�܉G,5q5"�VV�;\l�ن4��9,φDH]��P�� �R��?-ϝa̳ȸ�����V��k���~�7�D��}�Ό��?�����߸�IX���VY	ob��gze��Rr`D�NC�����͏4�Z<�> �g�%Xe���`f���#�ʈ�)�c���&��ޔ�}Γ�z�j9�3-��pY4΍�y�E��ס�t��^RgVh�Q/G��F. ţ��Y똚��"����v��t��	.j�,.��%`)���p�p���ʲ�u�dyF�'[Q�}'J�ޥ�5!j\Qrc�K��v�����	�REj���i��H����G�eX΍���݁�3�/�T�:�r~�,�7��R���e��ȭ0��B7W���ኢx.o �n�^V���� ��<��Xٖ��p�p�$��e,�]^#�l�k���P ��UR�I�����(ә�W�v���6�$#���Cp�� QvS3	1A�/�
�rtfs9X?�+��Eq���rE��l���ha5|���6]�Nˎ�,����%C^�M���#;�E_uҫ�ڋ�}���[�~�>$�x�'�dGr���e��®�ŵU҅�r#8J��S;01��ծ��?1��!��PQ':���Dٰ�!KѺ���ftge^M�)�f���ߒ�'�*��{m
��o��Z���a�T5�L�'~��^9(��#Wx8ȳ��!��P[���C~5F1�E�h�6BRR[T팣��Q�
����Rrz�G��%�bi�x���t����i}�`���:5���w����q3�x{h
 r}G2)4U֗��,���I)Zg&5��؝�׮��%t�6����4�;Z��V�g#2u 'R�H�NO�ީ��H��N��WYv@�lH
�������>�p�ŨI�~q$H ;�&IIDbe)9�x�@QMaµ�Lt�e�=�p�@�^�h9sF��^�n��_p`���!Q�rL�|>XA�O*t�����q��R	�D"�T����w��JB�K��PW/����q��W|Ǟ��y���:����p��rQ�1�p�X/:�sexPYJJ�7������T�{o젷�� �����d�a@X�"Z�,��_���5��`N�OG*���;����RR����#'#΅xI��1���C��r8�2�@�� ��+�����<��U=���2���$E�EA	}���	�V7�#�Ĭb0�f�+.�̩�wG�I<�����pq�PH�A׀u��ֈ�*zy?�>����u㪦U�6����waE�b��#�DX��I���g���!��x�����*�����o{���-w���������Mc�
�߆�T`�<Vt��R�ވ�D�<2�!�H��C�V)9+��&	���j*:����ޑ'���Tr���P{C�CRk1Hُ}Gpe�j�{���$.l78���{^���HGXCj_/�~��?>�'w: t
/9�xo�m���(��06����X�Dn�E��g��@$��iU�:�]�~�(��I�izz��>ˊr����[lRާ��D鷺ؖ�ƫ�\U/�.FbV�7�s>�f����,cׅW<��`��ƹc�QpP.0ˊrL8�5���G0n��LYg�.�;(E*"�Ҟp?׹�V���l��m5.�9@H9������kv�W�������*���V�u)6ѳ�qr�h[	�'�_d�0מ���u�*Ĕ^�}GJ��v��Kwb���Zԥ��\r�urn7dcgE7v*��O�/������|��|��o��~��je��<����c�
�R�X�W#|j�������&����G1l�c�r�dO�RإjXټ�c
�6� 6�l3X:~?��&�K��E�ƌbݱᥥ� L<�Ū��7T���<�X��Y(=�'�˚�89��!; �PK`4Fj�-C{�s����;��dQ��s�I�\�]1���-�Z����~� phxpW�,aSB�9!y.���2?F��/ḋ�Ԝh��<��%c���T�Y�ʗ���F������bs
�>1�b��4�]x�C�R�R	���J$	����:V�,�������"��z	7�>�O�ْ��J�!���?oA�Ϸc�ųV��E�[����0�a�����;];��@���H!��*�.,�
���%sۻ�[��]�+��D'���xE�Q������f�^�~�֭�?����f��t.�-];��qړ-�~�T��6���;5��FI #䃡:j�������~~�yw���4s`� g}/��rlܸQL�U�n�m�oh.
ݠa�����\a`8���H������7v%Li3���������U����;gޝ�`A��͙37�|3��y�MN:��> C_t[W�,<r��o�#�,j�@[��p�Զ���x}��F��ؖ�'�llOJ���z`�:
��������/��b�1�k���^:(%�(�wމcǎ�Z�B��?:�Ј����)�l����C�rb��硱�N~��d���Y*x���C�0�O���P����@�v�0lKˑ����E���$�g�%�E�g�9p�@��Č*����C�g?�6o����G��fa�	̸b/�7�i͌a[�.�'j�����I�E6�5�d��uHx=�#c=΍�=ˊ����+q��a�������w��W��_����UW��===3��Lx5�Ç˪�.�|a։_��W�~�zlڴ	������o��1�@��+p<:�ɰ��-����C�aj#Hƫі����zĴ�S�����Z���¸>)����,�7��W��oƉ��,�}�7�ݐ����ר߶m��I���O?��~�e׶�Y��W��������b�вQ�=�W��1I?N�����p��ch��Ese�T%*��.�� r���J�\��A��g�>3��efs��UG�**$�E*�=jq+����3`��I�G^��W���{�`����jۧ�S��,!?��Op���˗���ª�*�	&9F�������W��^�G�i�r
`xe��ѓ�zeKN�05�*�Ǫ#�����a
�(�s�ŒM��Wd�,���[F�᪶j
M5؎�
q�c���yM=�h��g-��F�R��~YY" $}}}��������i������ǽ�ދ�˗#��ʧ^�����F������'7�t:���ڥ)�>��+@������K�;\j0A���iG� �t�	f�((�V�+8�3�lb��Z����.��9��lB@-y��h�0*��$��/��N^b���A�S�b����oK���m��fvww��'��m޼y"-�!^OZ:ɠfm7�EZ�c"=w���ʔg�����fn<����������?�U��^���x��=Ԁ+������.�6� ���=Ś��.E{����Jr�/u2�@ngE/�x���_X���[������d����3p`�l.�ܐ�@_u0�'�E�W'��5M�=��l#x���")��.Y�;{d�=b�b�0^ӂ��s��zժU��v��I�r*L���6���QV�e��Q(��7P��&_��&D9sp<�+S@��P�}E�_WeØ;��5���5X��VX�1��k�=:00�36g��=��r�#S���2z�\�qÆx���H\�zL�
GM\�A_2���8Y�FZɋ�/�2}��ſF������VU	�<$�k����?����9��ʍ���S�ܷ�����{F��݋�I��!gCw�u{�O��L���'�>�@:n�|�ʾ�n���^Gx�1կP�כb�Qϣ
�o�l0��C�dy�	�֦�h�n4�xV�������u�[R�(��y�Gp>�2b�h8]����孧���TkSs|4�ZL��% �Q[APt���=
˗�q f��	��+J'�M�mz[��V�ns���A0CF&�C$H���7� K!�k�b����O�'�qi�%dk�&����S�8 HP;�!���c�" �	�~-��Gҕ�����q��Fs�Y,p�G�&V1R�]�=|��Ge@7�☗l�D>�&�H�`�sK��� /v�W�^�0�� �}��*�q���$H/�������G� ��[w�������B����l �(�G�������&��@�b�    IEND�B`�PK   J�X?��O�o  �o  /   images/ffe61187-e64a-4024-8cee-95dd034d2257.png -@ҿ�PNG

   IHDR   d   �   ��z   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  opIDATx��}`���ݽ&�ԛe˽�;lӻ�5���P�$$��z�!�)�1��ƽɲlKV�~����۽��tw�-������v�yS߼y��:���?����V���O�q�J=~��g
~F��1:8l�p�	�1�A~.��"8�� ��W��b�l���@���s3h������az?zz� �S�?���r��=�|��@e=֑#��!� 7/��j�����3���7�,zz�-���	�+pЫ��p���Ҥ�~�c�͢�ഡ���g�dE��I�7�~?�=���
�dQ���i�9�XY��o����&g���QD&@~푱���(�`�$&�.��긌�O%4<����ϴ���2]���/��h���0�=�Ֆ�ȴl�}=CI�cJ�3��6�	+������ޫ+����~W����YPS�"6�5�pwց�*�F��S��t��e|���VI ����XY|^�������g�}hh��>��|,�
��}0 IAB�P�$BN�vR�JP�]P��Q��>K*`�M`
-Ha��Gp�"r�2ɪ�}3�p�7�O�A��{�;.��,��(2km䢸`���b�	���Q" �o���Or�@�ߤ����z>�i�g��B}36�"!\��@��U#-T�15��%�CH��N��&�q4�wkJ����~s�#1���§W5¨,�M���@�f㳼��e^8�7\�0lLU��5�T���F8g���V����E�L��ϧ�a�����SjC,�ק���1VUd�&�{��	ɦ*�M*{^|N�>���=5.�}��T��Ќ�B�.���VH����7@�dO�P�n5�]�Y���9cݰPl�s�I�N�^	�y��3d�� ����ۀU&���<��� f��ŵb���\����b�"_�T�}���p�>A��gnY~ %&+��=���³V��ML|Ρ��}�GU�c��j%�=|T6�BiU)>�ϝc���-�@�;�ꏽ($QPg�)�7�>�^��Qn�g��Z�o����\p�;�6��(�� }�k~����� *��2�e��������Z�ʄØ+	�����g���{��E��c�2�c*��)�-W��A�}p�0�2HC�7@�/��&���f:T�>H,��Ud���c�
<6���}�^�d�FG/d�	����W$�~|�����Zdܺ*}i}�Ow�p|��/&\�����[���D5̝��������lcO��x�Y�>ϭ*wa���h#�q�@�e��<>��Y#��$*��[�����'�破Q�X<��2TRˑk��
�[�HV`j�~�5A��Ӳ=�G�z� h���ށ��;�f|��	2�6ݩ���u" �pq�l)4��! ��OH}Ы�{q��ע)3��H½���Y~P�gB"9.d���^D���4a��Q��u���U%PPsI)��a������AZ�(�I���EC 9F%��ټ�E�g$ꞟ��zGX1pS�8Be�^e8���w#{�!�l�a�7^��D���a��� \�%�J7�w�]�$c�_m�Fl�����ή2	����>w\i}5���'�Ҹg�܀>B�ۡ�c>��d7ͭM�&b�F1@�O��ᶩN4�;Ψ:��-m��V@�(pKN�����
�K{?��F�	B����27�B�lwGO��r�A�������&:�������bl�%C2=[m݄�g��'�ɲ���@vU$�Pw�N3M�U4��F~��$��Qj�CjV?~�'�h�&�/w��MBX+KDMi4���ê5(� #F�뮹|(*e��#�R�$���s��;���9�g�Yg�����~L/5�;+ެ�E=Q�).�O?\��hdX�o����_^i�����h����L����a_���)��K�n���ݑsF�/E�/lB��S;h�7��T�;p>*����o;"i�mP��+*�j���B��|عs/2"�8x�b,fHMM�:�[�&ޯ��������?*Z��0|�`N�����a���J��>En���N��6�U��0�G{���<�ѻ�/_W��Cv( {���wyF(A���� )k���dp%'ˋe����jQ����n�'$Ҋ<�TH�����RB���_��u�Lbl��*(�?���|d����Ñ��Px����W�����X������U�a���p�ݷ���'�ۊCF8�&@�	���*s���'���4����Em��^����:��Ҽ�V�A�`�­�֡�V.���Y������K��)\�%����kVc�-��<��o6^>�w�q�x��8-����$''�����M��$Z��=�E��y�^M�5t�4��H\ѳ�+�����Oq0g��sI5D���W�wz7�b��@��#�c9N"�W�8[S� �D&�cU��CB��P�Wz\ቂ�����&�=�ڹCE�'g	��n*JZ��EV�Fl��^�.��<HII�%K~��*��\�������l>]�5���~p�/Eb����s-�8A�P}2���N�S�i
��b_��8��
�\��;,���V�%h�]o�o�F3ģ���?�X��E��2F0>�ǫ*F4{��2@;�l"R���_��o㠰G�<�&�ڈ�3��f��,��d�F�4�l���#�N�1��b��Ǖ�r����l<[������0W���C�9hP8���8����k���A.:�<$z}���Dp5*���m��}t��w���j�#�����&QE����hxB���+S�`rl}G�þP$��N��;��I�GUP�A�x�����l�/cQ]L:͐WQ�GG��/���E{�p�8�A�O<:V����"|�r�k$��.D FP�D"+>�
7\G�ǟ~&$Tn�����⪶��#8TlQ4��=���87T�H�K.>���p���g��A	���D����n8k���H&py��
�p��)0{�P�);�M�����ol.���	���a�K�o����u>����U���<D�k�WUoC�����Xm��mHe?�>UpbL��?7�C��獛	ŵ��5Qƴ�����?
�`j	���&M8z,�"�qDY���e"��'Z� �VyME-�K��MLM��@;�*�=R��=QA�e���M?�,�^6��>�l��XZ����s)�"2�A��sƞ���?�qО9�$�j�r@���q�$5'
;e��:�D�I�d!9�tq`��U���r���D3���K�Ez%X~�]8�,���]��ӝMI�������x���� ��MK�M�ε ����½P�WFNqCg�D�煿@��F
���o�&?>�Z�4KJ�N�4Ձ�h'�FI28�/Ě,��#H8�$9�1ML:����&v"�dW�D+aA1z�B"�\�R�ϐj����\���b���_	K���x5�H�A@ܠ2�a�Ep���Pଆ)	bM�Y��|l����$�� r���@��?]�1S720(��?��5�s��i{�������i��}�=��Ͽo?���I>:����?��&�i��2$����%�����R1��	�6%|`��M�q6�P<ƍ�ښ�t��d����O��专�_�_@��J�H!DBD4d(m�uL Hڧ+�v"��d����=��^wh'�S|YW)�a�ps�f� V�UBo���־���J�'���A�4�N��~���bI�^�!XYm:G-^�np+�����E� ��&�G��,Q�4�e�dM>/<_Q#�q1ɒa@ب�1f�K;e����nuX��,��#�0��0'��`�bH����&�E��
���u��(0���h��c�Ǘ���	>��򬲁d�ǲ:�/���5�Ϛϐ�D�+v�{�Wv5�~������!;�C�֭ �,pY(߁����,����`��<d{�.�!�s+�B�dUg�`B�o�_�$N=c�[Pz���A%�A`a�E��Ų:p�p�D��!�aGI�2R3��q���-w��S����H>l:���L��	:��0؎��4hlD%������tn��.��N��&g�,͇�Ź�x^�#
�#�U5H��lF�*�\�:_��h�����#`_y��GɌO���x(#��5,=�[sGL��yy}uk���@�%��	��a���p"�ݸ������+�y������G����	���t�QĐ�J"F��&]b0���t�F=��Qn�=t�I>��g���Z�4��[���{�&�C")5���˺��"to��� �>��{�WM=���xrВb��	O���ѳ��蠜,~�9Pd+�e����s�Hx��[�
^�?o�g"R�1Brq��火���n]�mr�}Ӡ��:Lv����J(�)�8b�YӠ�����	�)i)P-�x���0Mh~S��qEzdp� 蓀m���6�hn��%@Ecm��P߲�)P[Yퟦ��48�����T�p܎��w��A�?��O+=��[��Ы�k��^��Eވ���'�?M�w6|�G)!����/�DF3,ݻ��hq{�QC7�9���)4;������χ��۠��+�u��O�������Q�ז��h��Q\��_�X��h �;��б�6x|��;��p ��?ݷ�G��#�U����$�Sƻ�|�I����&N���S�(2�q2� @QeQ^]D�k�E} ����	�W��2ma���nW��	�G�n�'�~?�Ǳs����<џ�7��O�B3)2��N	�5A�qb_j|�.R��c&�gA�)z,���&�R�+[��>.8e�'�(%�#��Q�M^��#4�@��_�z��S"pU����t��t���A�D�������N�3�_�8xV�7YJ�=�s�ֱ�d���w4�?,�5�r�1r�[}�����	e\$:�9��ף�36.
Q��q�4y�Y��	I�+����/C����H�;�k�����D�	*��&I�����=���*F������v��^��j��R00�������n��<��pEl3)!NA��F�;њs���ʒ�/���p.��Ɨ�C\�\v�Y�c'�>�%�+)s3�;Y��gE���î�"FWھ?��,��cgK*q�r�'#O����������F�W�k���
��.a�Z<���;$�Q�Jf�WEٽ*�h�]d��^�>p,<2�rش�4�|������9W�}?�;Kr[���dr-
54Ei玉�O/�{ecu�}$���wa,��N�mMu�:��Ip�Q���_��o�a�*��/ �?&��z3T���?��t�Ȳ�S�Z�r����ϛiB�/@Ѹ(��h�#� te,+(��AY!|.��Kђc;"��נ���׆�߹�R�{��t��#+�8X��c�YjS��׌��9���:��5.�G���y�0��}��1B8<�s�(����҈�C�_8p�;Cen��fZ�k��&�n��*u�fԣ�-L�V�8�rZ�\KI��j�����ֽC��8Ś���j_�!�^�J���63��GH��b$q��ə�@����G~�>���"��zb: �ÿ����x��f(�v��xTB��>�� P:�Q���;��楂ݨ��Jl;Ú��M5\iw�H�PTl)���4qNo������'��&ua"������O�1�4����W�R�{$��z3��Zc{$��;UByC����_�Z�^�!R��HKi���a�8}Ѽg��isS�O�=�;�����\�fw���+5c!\w�F��,chىh3��Ɵ$��+���#��V��N�9Yt3рh!�k��R��� bг���Y�qM��M���[K<.�'m�BZ:���>�`D� >2��H�[V�Mլ��	Q!�]gE$^W���V����7W}И&�#A���T!��צE�5 �8�m9�pF�K7�nm�}?�U�T�Y"k��0Ev���V��;P�Oy�xl�=~�'I�eW6�E+�@�kp��� 5�<�?��"q�~�/�p��LY�8���a�y��!^ji�!����>q����D!�T�P-Cz��Hד�¾=y�1���;�.�`��e4�ğ�A��gZk����M��K��oM�(<i�U�( pJ��[�<r=��$QeCu �Ac��\�W8��i�{jjj���D�L���Q!.6���H)�~���6bq��E���\,|�#�!��ґ�F�^F��j*p`���L�M�N��J����!�|�U>��G�?Z,�u@t�?{�,(���ꗘ��w��&����
Y	��i�O3���������<n���s�����Cae+Az�l'r���(�qDuW�eQ��N<���f�~޿E?��Wь���Zp��0b��V+��1 )%���������Z]��.�eI�|�2XlX��߇�Qt�x���8Y�� dG���DN("J����l�R���@�VE豬H���+F{��� ����{K��,)-��q�h�V+477C^^^��s��U4-���a����F=������?ڣ�;k�IPX[c�PLaM���lHg��&���u�_C
B6�$3w:�?�i����3�����B�dG%���V7ќ|t+kr�̡ཌྷ��$
���%d1���@G�������>��l4h�X�!�}��v0�D33v3c��h�����w�DäkR�R>�q5e#F�A����r�r��-#^����so�/����I�j�@R*�3hLmST�z|�s������O��p)�.� ���;��]�u_�n0�$&|��0ۚ� E}#Nɢ"�h�|�)/���\}���x�RRt�f������x��F����������zgL�X�>���&A�,y����~� Uop0�`�-o�����d�7O���)����lE�"�u��>�t�zm�pO����d�}��B�+K,��D%�qg�;�D��Mu0/>ŇX<:A�DJV�2�᪖}��^`�GUO�������6�5�o(���dUD����o�:@i?$��EVO���T�S�6=��RA�{���	�f�ϩ��XO�m@8#ܥ�7Tz���.���(16'p=��~]_��eɦ�+caV���ld���Z$ưZ�w��m~�,/ k\X�P��6��hK�v	)U�
a��תD$�~� 3TGsj;�/8v����e!���vl�/
�Lټ����|ދ��7���J[7$	��|�e�G]P�_�	�e&��M 7^C��g[n��GS�,���>Z�#2���N�C�(F��U[��W���ZE�ar��U�b����͋�J���HEJ��[�#������K!r�,�yG31{8��n1���w�_�+49��9b.��	q�����z:�Z$����q�i��,�Ӻp3�9�)fO<�꒮�\��]��P�0|mVu�^V(�(9 ��\�����C���-������BjzZ�*>�@�F��s���|"'���
�����́�hi@���jeti,e�}��������FmC_����				PYYɿG
�P�dРA`Z�+](z� tQ��ZH��B3�59�}��>əPUUŉ����z�����п^d��-��� *��2��D�$��P�O:�<7�-�x���ƗF���CEy�; i(���%P���zp����^qL���o��C#�2�%
Z,��g�^f�5��kFD�Dv���]����lXͨ�o>�T�q\�qr�$��|�!�u�PU_ó��$�Y�x�7>S@ԇ�Q!_�y��L�d䎚,�Ů�@�.h�H3�$�tN����fbY}T�����w`G��4X������4i�9�&����9:Q�>)u�9��7�������!Ȱ&��P7����q��[�-ű(���v:[p �]XW�m�
*Ø�*_����;�*�Ѕ\��9ݚ7�e�;���,-'kfp34&��F����NEYo��g:#z��e��XQ��E`��	i��lk���)���~ˢ�N����D"�\v��&p�+�Ԗv]a~�=�Ó�K��#�]U��<9qG8|Y���ͮ��
�V|;��B�,��jɥŲȃ�eڶG{�H�x5�����:� �/�E�Úo��Q}��~Z�W���W&	��"o�~Q8�^I�j�N3תŲ֑>N�4���%{A'�h@sOR6�)� b��Q�aM�7���_��^���*��m<� @1u��i����}�"g��|K��g�h�ꄻT��ʛ������M��j���)-� ?��$��.���,H�#d[�l��ۯ�s*�i��W�kmŚ�g�@�����@������p��h���߼�M�����L�3�h��벪^ *�E�(^����*�A_$��H�5�uPJK���~4S�\	�8��i_)W{����A��9R�3*T}a��y���N<�V�Lk�d�0��1��bF�z�|��׭�VkyY��e1p�]�t9[^���C �n:�B�ڗ��d�d���z��a ��x���3`|�`ȩ9���m��x�Oܔ�	��CA��@����I��ՠ�܁��cP����Tmo��6~�	$)C�)Lh�P��
V�W�>�����Bx?�#�,��ƒ�~@K���>o���d�WR�6��b!"��8z����êO���
�A�� �͝��S,Z&uW�PP�jk��Y/kӱ4ge@�M��6�^qj�� S�|Jն���B[{h�!"�o��NZ'��a��O�Ao������9B��Y�p��&kV$c��)0ޔ��*��F�z��i�X�t���\���W ����Z�G;A��'_I�X��ʏy ~��F�RSz�i������:8'C��I�,0����c�an|J��5�����ʄg��r=�3	i����x|�(K�%oT�T������Ñ� �	�(�k}���"a�8r��_`�޵�0KQu)U�����N�M�ߥ�� |�?w��~)���DK�L�.%���T��&A�.p�����c�*�7�LL�q'rIg�$�$�^��Ce�<�VD4n*&��s���(���-|ݛ(T��}�r��w���1�ť���k���A��$����x�E�F*W父�-*�Д�Yj�v蕀��֛R�W���z��\�hrۏ��Ҷ]M��iP�d03��ZE�,7XkUH�5vTR�HH�O�eMs�J6,K��}5��3-K�]�\���@��'=�9��53�����ǧ T����Z,�p�b0^�,��͞=�[��ZZA:�9#N�����o�ȿ<=�&R,k�K��!�����%:<ͫ��d�Ɍ,/�����?��Hj�[pI�S>r�}߾ڪ
�?t�Q^��
n3�o���f���x��"�����3�rU���v������F}���(� kNIfM�
W#�x�G^�&%"©ԑ=Q�#Í=�)���#��"�P������3P|��/iu/t���'�$}�u�9E�<~��c�C"�ߵ��l���M����*_b� nKg�w�=�{����1m�I:��yYv-�xQRD�to��B+��w�e9Ƕ�� ��{�lWڼ��f{��6ӱ#xd�}�,A�4���	�S�	^(˷N���s.u��@e��1p��S��� /�,��Ei�� ���?�	��H��B��'H��Y���A~B�{CM>l�/�y��c�]z'4fD	"�͂o�Bz��C\`0�32�Y���s��k1�!R߯)W�)*��[Y����Q$RRb�u�� N��T!lUR����2�=f����,	itU�x�X�ɼFth�H�H���qԠr�7�B�h 2,G\�A�t��oEX"��Y�Id�z�"/51aa�m�ԫ*sЉ)��M�?���G��&"
-��_L����O�D�*�����z�%��mܪ�[�(}&5Se߇Ĳ6"�J)�\}���u� H�Q(�e��z��i������/ ��"¥�q9S��_B�����FtJ%��ԙ�:ѩ(Ih���\XN;���tgI�r�"z ��k�����8D\~�G{�L�p���kaF� �H��f&�6D��Dq�r!ʻQ�]!�>@"WUW�ּ���A��/����v�c�h۾N�O�nF�Dفz�r�!t3��mޖ�T����Ak����s��q����`dЬ�H+!;	�@��R��!9��������Q>�8�HY7Wi<<T?b:���o���	DI�V%o�_?�8Ύx\�$��W��	gզ�(z@Z�u�T�M���
�m����>}औL�gn(�-�(V%(���9t���D\vJϤ��n2 Gg�j[=ז���!<����%X�`d� ȯ*��Gg_�7~n�w��$�����u��Ⱥ/�E���$��u$�b�ŭ?���90{�$8��D(���K����F��XT�֗�[<Ӊ�E�Y;p3\cתQu%� Jg o��0A]V
�I=ȸ�`�cR�Hi�ym�������[�����Ǟߕ����'�m��!����M0�2�Z8,Ԁ�t��g�����J0���Y��/JCi��,�� `4@������pZ�KƉ<Qc�_�Ѯ@�P�&z��I�Y��!ǰ7]�t��U�C�-f/�ߞ���}�{�W�@����7->���xE�5kւ���9�p��>ْUc��22	<診���.�h�����0Y0�$NKN��x�阗��hթy"���I�]�$�'�En��X*�JLL�~������#�_�Q�((/��c�B�lB� RS`��q��Tղ��I!�n���7(o�^JC�A/�Fb/����Sx4BU�>�<6%ů�lN��\�r{�0Xok���r���i���57�s��I�����[��g���E��L+��XW�~�2b:T֖�Z�ڈAbHF�6	u�����;i�}�x(u��K�?�ha�5�B��
_�o��5y����f�p^������ږ��bY���k�렬����(�H!�DE�/�����4+
����m��B��6T���^�R�޶j!';%,L�����p.O�얍�X�r��ؖ�rm��(aSs!��Vr�A��2�U����lv�� ��L�~�$-�����,�4D�e��g`GCs�+�˰#��%N~����!
�|~�����L8�/�u^.�d����#�7����]h��(�=D��Vm�V�����ے�Z��/?E�`�!�X�#c m.��GLц`��#�<,��(��r~�⻑r�ZNB�OU��{��0Û}uAR�Ϻ
�>G�GK��Hɑ�v�� a�	D!iۑ�7�qG�X�Ze�E7�e�U!1�F�6��Q�ۓ%�[R"����xP�d-#ٚn���(C2^���8��Sa���P�TFd�ԸDx����2x5k�l�0	׽@r�r��Ғ qG�ŏ�K�N+��<䒵��b�����������H*5�JzB�쳠A� � lF3��6�_�S�L�g�}e�� �o9�:�o(�L�P��@���A���� Q֘�o���;�ċ��C��@����#�q���8q�y"ݎ���ZZ��m0�"�k	#D��{���1��� ���� �1	��-�q��m��������Й��%�����{�RM�"7%��<���j^�!9!ds|����8��&Z�3�BU���"�0f�Z@�ά#��nH�w�҈~�6I2\�o:*��h�#���dS���ǡ��C��ʦ�2���!l)ʁD45�>���3zee_�Z4��A�dn�c�C^�=�&<9���
Vs`�V���P�:ѧ�&���h��k!��z{���a��Ŀ�O�.5��bY�k�S>j��S�(>�j��6��^\W/Ք���8Mj]˝̞�%��AN�z�<�+�PS[
Yæ�6~�5��n� ^h@o�5�7�ldK�:@�`oh�)�?�ᆑ_F��T�m��q�HJ�!
�����*�[S ���:�d��![=8z�o��R�{�ύ��5�Gx��N[�{�#�$Р��Z,+j�\4��t���a���Є>�+�I����~�s7�p��S�Jk���À����~�=%��t{�.4Kr���qr8_�z�8L�0�d3�䘬�����!�h��g_��/�i�
Б�SQb���k!=d
��K�8%_rֲә�
���I�|$�%���B4wq�k0���q�`���6-���7]y`;��%@ay!<���S�����j��w[I.l����-�F�N��p���!�[vt���$��#�?f$I"~$^}�ǡ��:>��N3���~m���jQaoDT�*���b��q�p��Oj��Ъ;�
�X��0Ā񂨥��j'������,Y�����H1az\��զ��e�+&��@-H�k��a���/xp�Lk��W�+q;���%�ǲ�	d���q	�d;q�_T�.��4�(����a�@bd�b���TL� �� :�$�j�-��EJ���}��ы|.�|=������9$&�`Z|Qr��i�)�a4�<���|�"�em*���wah�{��&x�/!^�	B@=�N��Ę���0⎈���� 9ā��d��� ���GU�l�{^*B�������fz�q|��Fƶ��:�d�*��2��k�� 	�[f_�'^���[g-�7�-��##��h��(��[�vt��嗾�1:s]�3�Ųތ%���0S�V��J��j�ݭ�����f�h/x@�Z�АB�SDb�(H����zO��Y�i�����+�Q}r%�]�L���\nXbL�@>�_��8Fp:ܜPԖ8�KA�1�W� �3�]
�#.2Y����b�SI�3%�6��#QD����_
��C�,l|�jt��촃�__�\ҹpŤ�|:uKQ.�;���'�@�N:ÇD�XL\d:bb����8�d6p}C���AXp�{��S�g��3n�?��g��kR��+2�c ld��uv�:u4����~O����~��
-L��D��ZXE���(tJk�់_�,+U��u����P4��C<��'� ��8�5� 11������>�lX��b��\|>����'��p��"�_�8#��������D�e!�@��-}�q�<o)L�w:@�捶O@�G�[�����T\���!��;�9T��g�l���-&�^�kDh��
&h<0�ɆX0�{�G��5|*���Q�X�o����E*w}z�l4�I�'��R4��g� ��	eu�]n`LdC�E�)K�����ne����22Y�o���(̐�f.�U�oc��@I�r!Jc��ѫE-`�ʺu�\�����ҽ�!3!�ω�uQ�@����!���"�n�:1j��脢�ta��e� 2Qg1͂��p@���w�$i��z��R�A�%^\�Mp��+`����ܲO�ˁ��("H\9Њ"L�m���r����p�BD"�ߥa���~�h�����G��}�Jhvt����ˊV�'R2 M�o][6^Z�	��[�T���Q�YQ4�)hH[b�@���(�z��1����J�p�t�zq4;q  �/�9*�7B3�fbќa5�+��yY�$#;=I�*iP"~'Χ:[�`�[4*���zVc��W�+�v��N
�������oF.p3�]MF)PƜ�	�}u�?T�lW^ }�B����E�:_�}�C7`rl$�_ş��z�c1>�&��^��>&��\��4�=7>%�bY�WX�h�ѧ�3D0y�>c7c�Ez�r""��ڿL���������4����@M�l�^=�
�?_d��}�0�y,���\��(�Zx��$H�����.���E�c��6*�6�ٗ��hY|qr�Wå�#���}I�6��yy��Ě>hL1[�������s���ُ2�K�w�<\t�xLK���%�H\Lu����ט�δq�����τRڟMD��p}��{A�(ՠ+q*:���8���v��o?"=�q�̋*���mS�K,70a��Z�ƫ*��7ZfX��~�lcm����-@��������ִ�#���ΊK�2�a��Q����ƴ'ӱ��G(y�Ũ��*\�wm�[�͂��}	e���a��X@F'�?U�F��pj��2_�˝o�U-���y���i3P�� j!dMB���"$B�E��� b���x���6@bR:\5�t����)���(��n�_�׋Re)��N	b'���*D�{M�4�^w�/���c��'�����̈o��f[C���o�����#Qƃ��S��ޕ{Yk���~�:��ǎ���(G⨟�o:6��Ecu�xM�����D&�}A�K��t��8��9UO��+m��f����RF�Yl�Y�Q�p�Zp��������w���w�D!��.K�s?>�JdnC�ވo?%��	i���Gh���k�o�߸����?��o�<WK{� �O5����l��@Z�;�yH�G )k�ь��B�Z����uB�d��9���m������F����;�$W��v���U�`M*7��u�1p4>�pg`,�k�s��a�Ixx1_cx����e�f��ݎH#o�<o��^:��K�{oYTR��c�Q�{]���_�A$�9�E0����@h������-�v��c�>��,A����
b[r�1����	R��J�/�^��?�9���RT�F��E�J�J'&�����c>9 ^���H�u�|�&�d_k.��<o�Q����)ZҠ�����h�����X�� "@�4���hL�lg��I��*�O�\��i�;�s���\w��n M���^��>?.�s�V�+�':�_m����I�(��;�?C��ޞ����9��`,���a�Q�G.)m>��X ����u��Vŷ�Z�l}��ߙ�M���H����F�(�5U2�	im�R�e�q6�[���x�
p��O��e��,�4�K����i���mus�,(~�/�B����]�o�&t�Z"�e1zc"H����Br��anCS�yxa�B�#�b����ke�E���d}�q*���[[��uK�c-���M\��K&tw���l0­�`�)��Y��tm���
�R��;��(���{�ιdU�򶌁_�RY4h�9v���}&�QY���8�2��yW��%h�ъ*w$��@m��	B�-G )�1w�Vb4@��pg��[p[ڀ�׫�/D��&�F��<s�n���%�����+���[دeFA����B��_���l�y�M,�@��Ef���9ẹW�)C���:�yR��������p��#�?�8.|���r�����2�����]�R��1�.	QWkN���ݺ.͠�hr8%���@U	�?n&Kφ�YC`���G7A�_���U��8$\J����F��Z$�#�Dj%l{�A`�ă��'7˾�D-�u�Ą���@a;r��MPgo���WV����ˢ{ g���2D�V��@�E�����YPe�)+�_��"���w��Ef+m���C�x�;
��=g��ν�9@��,��<-.�}#�Q��͖̀��j��\��J7�4��_UAk�@�b /z�1&�ڏy��т�R���w-�ڛ�8^@bka������B�/m%��ɤ
4ދ��D4�<������'_ k�w@>rȩcO���P�uG:i+PU> �d��+�r���~�!������F��
�z��?O��fW%�Nw*����h��'͇��)0w�xo�w�|!�	2V�E�s$.��R���8����K8���.�e��C&�9cN���#��m�awI���#d!".�	5�\dUWBIsJ�.X9���R;`{��i��wۗk� 9n0����	�����"�҃��>�S��x� M��O�/I�OCGp�_c8N�X�59���@[�@���B��t--C�KH	L�c;�q�<�Ar�s�󠲹�+��hr��7C��w��N~ބ�$*F��.h�1�<�X+��Maa"Dx��MA=cn�� �iC�%���Π$����G�ʗW}%�e��0�3%�Y���q8eb{\��`b"\�:-�>��]أZ�]߶Q;�bM�R�"��e���tދs�SU>51aRw!��#�<_xю���*��=@H��z���[v�y(e.w�J�E�@C�?x���F}���yP�aB-��Fֺ����(/�(��(���]�����o�}!ħ2��mR/~EJ�p(�E�� 	@;�I��M�V�P+�{�Y�螙�c-/�1*O(�>|"��z8D��n���A����I*��?n�g� �!�T�֊b�L�FN�f��F#w<A�r�`�KQ���:NUكa�N�53/��5h�ȋ+?���C]��������}��~B�$AJB"�x�\x}��=�� �������Y�t:N��WQ�̌�d�⤭����C@���8m �O��J|R��0w�d�Xǁ�z�YY�&��!�g��I]��A˥c�4�<��}$U��6䭚C��m�5�b�[*���cY-��`f���R�����rz�8�*=9M�!i}ᥕ�w���BYC,C3�vD�?wX|�.�q\������U� ��v�m,_[�.I*Vdu�˦/hߵo��^�U�6��,�Ԭ�=O�xϫU/���J;�
,���.�@���cm�%D��-x�@�W��?D���'!�~t������B�e���xQD�Kʀ?Ͻb���H���x8^�e�sf|
�m楰�� ޤ��y�2b�,=�B��a��̱	-��[���a/���1�u�ׇ��
H�����cf��"���>�����ᲃ��Z��?��jri�h��D^�=Yз`)f�ΖL!�L�;5�RJ��hf�֔�3̎��q�|���?�)���P�[��p�:��FnR���'�5�[�D4�Q�]����XU� ��|bؖ���l�2ڨ�'�9�,����dUy����S��GN�I͑��
3�N�kBN5�#����Y�k��'>�5*p�����	 e���>��x!�f�a�C����>��uhH=A����gNY~ �,V�S�{D&��g��=��{Ρ�N�xT��11�W)�U�S�y�K��a�A��,���O�����o O����p����'	��11�9���ʹ]+�H�{L�P����6�A�Q���<�B&)��`�d���iQ�n�K��)9�w�}��A�^6�S�y�O/��&-��`�[U������F&<�㰵M���H��#�@yS-�P�p�e�������[����K�B�%�p7?!�A�*�E��C�^�"k^P�x	��NE~P�2!����&��؋����/���� ~E���7*��N>�d�z�����_�Ob�u�E �VB�v`�z��Tz���
��$�%J��1���F�5��n����ūPd�/}�sǕ�Ws�7AH��DzU#'��bCR��;����#`���P�h������l�y_(O���J1*�l��ʋ�Ж�Q%���1Q2$��t�&w��'��~�
(L�@�(�gr+�xEk����z�̻^]MS�AV�����@�����e��M�/��;��6t�px�^7����ᮀ�jDvU��ǲ�ر<G��������B�,���x~r�6��/i���}���#��_c�$���C�Ĳ�
1��*[�k��p�у���AD����!�X�ǲ�"S̱�� ��	Mְe����2M��e%H ]h0),c�Ж;�>�xUŸ��ז�t����'��+J:��U�Y0)6�������[���RՉ������rE��m���ώOyݦ�_Ҵl(� �)��X������Nsga��L�o+�:���%_��s�K�3v���=�O� �a�K�o��.t'~���_��ɪ��WQ����p��&0q/�SU��-���L�>ź������mˍ#��'g��SN��J�P���M[�r"�/�cL<O��~�+Bs��T6T����z��oB*_�e����>E8�r*��C5}'�n$�����2M�c����NE��O�ͻ`���m���$�Ped ��TcV[O���z�D[3���`#�~{�y��Ew@.��w{~��w��x�:�"�©g��*i�b�5	b���
�3��;Uᦝߞ[�	,ܶ|nW�؟y�O��.���>����L��+Oy�7�BaM_���.���!���ֲ�3v�<��y5��j楬X���M�c���($�ϵEYh�0� ����p�	'���x*�k�+��w���|J;"	��Ms.���^'d���|��G���AA�H����0 %������]p\�������|�g�h��w���C����6��=�`g��-/#"�Wډt��SyA�/�:�:xc�bx�珺ŷ!��fYS��V|��3H�.G"��w����!)U��CPF����#i9�fˢ���OD ��?�TZ�$j{��Zu�#�,$g�#F�W��W�)g��z�z�rD���v��[�~(ή�r���`�swp]t��I����^r���c�jT!������"�Q��|�F�n�]�d5���"�(o�M��[-�i�ϓ^�"@�e�FJ��T&�҄|��VN�O���������IK*y��a2C�3Y���N+���j��&��\�*$!����`=��i�N�1�\�E����1���$��КuUi���gH\���^�������W�Hs�%Y2�k���i�']�)��<�� �ƒ�XV�����B�Q������3�JQ2�,��!�HE��>��g��5���qk�hi�#���Ӈ��W���s���-�0�^����
3FNF}d���gU�"1�y��Ho�)w� �u4A�(*��*,�.����Ew�D����������@���4��S�5$pYV��h�U�٣g���KQ7,߻>�m_�Pq���;u�/-���]2�,���^����Z�D^k�V�&}��F3t+D�e�]��\��ˋ|��yT�E�G�����[�t�<x�y)�<�C���z�O�ˡ]�ӯA�̓�-yʩ@M��LB�Y����Q�]ۑ#��-p:�5��=�`T'r(�7��P�	VJr ���X���4�5��\�B���Z�#�0��K�L&�\<�TxEQ z�+f��E����K��_�����8N?a�̓g\�hg���̼���EXG˳I�g�#G�Zᦓ/������F���kMJ��lF�n�Bi3�m��(
��֏+^�?�uԲ�q��8�� �CD���Cq�
Q�?��_(����YȈo��&�����J��W�2��F�y�{2�4x,���]�uh�]�������*��bY�3�RTtj���-�4�R��d�)�n��q�����[�;��hӠ�ڇ>í?	�]� ,��_p���hկy�v�p	m�l�D���,�"/���F���'΅Oo�'<��˰6ok��r���⒨���C!�pg�~WO���b(��<�y+VO<;1�Y��$~���C6@ef�s�:�?��m9�}��085�l}�=���GaS�^��ZX	>a�xx�ڿ��p@�x��?s�7�IL��~�%�w��E}|����_T�@8')��W���;��h��������H���(�oM-��*a�7$���j�ϝ>Pҧ�%<�Ccuۈ/W���ڷ��W��c+:L�=���ܯx����۟����MK���ԁ'��Ac��+a'�_NT�}Rx���YP,��r7ö��!���O���'.���Q�8�� #�O���X���wd^}�xW��K�ߝDm�N���Vb� W�اz7h)�TCEg(�hf\�QY�k��bR߂���_T���+Kx1�Dt�N5��R��́Ǵ(���u_���7��~N2�;�3P?�MpB� �=�ħr�po�!�D�c�R�]�3��mU�qڤ�A5A͜D"�T,{��D��ص�v�X���������?F0�]�r�ɓŇLBP� 
�Q��1/iC�OGGp��@Jl<�û���/��/w�`��5�����1��j�ZL�&{3,ݾ����͏qn����?�b�a�'/��=�	�����]�����p�aH�۩xW���?��i;Ol�JF�q��憇�Q�1���!��`������8A�*p;����B�1n&����cH�@z�kP�uGy&*�/n~�����h!�㹾�4~s��p���ܸ=uK�B�)���=��/��+�;?~l�f�i�jX���A1Hf��G����'J7� ��t�i�@�e�a���"�� �����S�R.�������9��Q`lL��]8�]����u�F��g����}l=�(��+��~{���1�#0[hO
���7����mPX~���a����mSmRJ��
��;�\U���S������}>�%m7����%>��>����IN��ɑR��g����U�Z\�XD����/�/����ޏ���H��ar�h���g�o���\�f�>	>�韐���N��@�_=��S�l�28�⌔5%�e'e��S��J�^��"(o�bb׿�4�[�\�>rEy��dhv6w��3���:o����j{Ĳ�z#���^��p,�ԩ�lB2LɄ[�� ?��]�^r7G,ͯ�����f&����p�+y�.�[䗐)�p�28�廡���-?n<�|��\���`;ꘕ�qB�Cn�E���ґ��]�Xӈ�W?�{�UGNM�6��p�ؙp"�QS�H�{	� �w�{��C�����w������z+�%y����[��(�6��6�m��@\�-3��]	/95�վiH2z>��Q!�d�62+��AK$..=��3��BQ�}�r/l"#��x�r�r����w��S��O4�z�eHL��"=��n܃&�.��3�6�h�k�aK�渓ٛ���P��a&�h�hg���hL;��;E��+����&;i^�#��kBD��J_�Z���;x=m��}��aS.�f�$z(t?��0���A�0���ݶ۬��&������y�f�ݯ¬gn�]��SE
�GL����f�.7Z��5")#��x))� �HDL
�������l��0x��?�D��X����8�H왣�����k���`h��B�Q�`��o��䓭?���M0������Ϲ�bw��89��L�K�ZA�����l|H��o!E'_�������\�W_���磈I��`ְy�E;Wv�jANJG%~'*g�����yP}ڼ<-k D��Ϫ�khS��
�VN�ہ��<j��v4 6 Qhn�4����}(�:ܵ��t:�C��oػ��b܈g�	n��w��xDB1�ȭ(�fA؊��PD��zG��׾\���[�mbgX���������QP�=��{A�uaH��#����2d<M?�l��e�����$���r�=7dHE"��9��'�K�>�K(r�g�P���rm>��2��f� ���B���d�;*B񔬪O���;��X�J遑���z3��Zc{$
"nK(o��K"���"���s"�����d|�ˏ������&+	I���"�Z���襡��qIP�w��%�0^���r��� E~���&K�����	¯Q����Fm�Ҁ�L8����pf�fR��S�-��F�{��B:�?8�o"_c�'g��_� {�c%�m%g�u�xM�A��$�����bU� �"	Ǡ(�܇�^�9�����%.�K@�k���<!.���_a.�:���hj��uɈp���Y�a�n��.pS�|�fW��%�JPD�L�5˾�uh(�Y�C½ ���zLZ���4[����ٞ$�y,+�$��i4yI�>��]�1�i��X��D��e8�U�ó�s����n�J�_��[t|5/ZWWͺ^��^4���24w)��vg���M�ͧo�ؾ�o@s�S�����9g�Dx��x���$�܀.W�*Ų�!�`:%�hډ?�������:��*���{o����WX$	VIT$VE��V0��kx�OYWAE�
��	3�r�!͐&�t�����힞��a�}�������U�:��9UNm�zmq��!Z��מ��W�X�V�y}w��-���J�%����҈n���?�ǧU5Ț�CۃZ��@����4�ۃwr��'�H��j5�.V�����J˙=��mRB
���X�p�i�p����HCs�x�-Ըn#y�?���r�e��"�y����#t�+�Q-�����7�X���k�|� �V�˪��s���^Щ�}��J<���\�/?�"���\��Ѵ�&I
~ⶡT��q59n|��/n�ﻼ��Ԑ���;
����^���gz�)(_�1�u���Nۥ?���/̥6��ҭo�55<�*�r��ך�s����8%�@�i���h��B�o��nq �sҖнzJ�ǱW�l�N�r� �-L��ǵs~����osdcQVֶ�s��zQC�5n�A6�:�e�Ay[��2_]L��;�3K�[��h%_�D�"��J��P�_��x�$�5[�5-Yf�K�!`!L�SW&=���^_>CM/~�� �_Á	�.N�<�z��u$;�3�)���,�a�l<�G����6�Fӂ��Z%#ːZ`llqHV��^�,l�r�Fy>�|���@V��n ���	�6q�<+1O#�F8�9l�&2B-~ ��c�ð�RU�-D�/+o�1��#]�̂دUahP7kV[��a7����-.�-`a�>��9A�@��j��()Р�ff���Ec��:_ۆo�6�x �j2D��*3�PEv���e��4�BG�[�@c��6�!䊥:F�������$C�L��U��t�DJ�X|U��;F��+�Y\���B�q#�Ζ�LJ�@ʒm��m�=�޺/�8#-R  <���c�*5vN�����X1�V䆊K�4$��̫ߣ�A��r�S���0�}��o�>>� 7 !�*�6�A;A��@L�+Qްc�\FSM�}G�h@�[H��ւ����$;个%�ޠ�s�J ��Z �0����KӇM�m��#R*��ߓw�� ������0/���[�<��T���HL�_hO(Y������*��NE��,��;�z݃���^��b�
�����P-�����`�{N�7W}
u����h�����s ���A��ؐ�<�#y��[�C���=���@�&&jE�0�P�_��(�3s
�^~�I�w��U�g��#�8=���缞eum�_��vVp0¡(�5���ڏ��Z��V���m��)�b[�O�0�xi���a��פ.;���e3�YjC)��=�MX�O�|t��[���������kgJ�����Dȣ<+5"6.���;��>p<��g��5BFWuO�#�� !��q�.v�6FFv}����0Ya����n�L���z��{0��;~ܡg|�m��^g�����$��-;J��U�y_LY���I()�1>�7�yz��8il�<G���`�rF.�zpcV�d�:�;8��٤��]�77m'���&�O�PF�'�f���L��8~x��bԂ�ߨ9%c�r}��]�n�*��CF���z��*�&�	�#�l�V���1ӵ"ݿ6VQ����)?��T���ke�f9�2��*�������~W�>������
ĳШ82��z�V��p�|�J=�5*a�(s��X����h͎t�E���<���r�s��+��Yf�v;UGu[,��B@ۨ���h,��*�=�vE�N�L�f�]ɺ涬��N��{��W����Vf�P�����c�x�ڕψ�]�Z�3xx�d����˺z5�1��J��F��D�u ��oL���� ���%\CR0��[���ƶƤ%�h��4SI��0Z�:Y�Fe[�?F�Ι�ZK�Le�Xx)pt�^�V�ӣ�=E��=�^��_f"�U�K��y�����LD�W� %�,h���?|����m��h���s��s������N�7�%���5_�|v7gu]��5��OӰ[��彄'�@B%�ʍ9-b�]�q(LC�ܯ��%�a!�*�/Cj��^o��^�0|��Y`W�資�&eրv��c��KcO{	�w�-m�~b�[P�KL�J��ʠ7�`�*�T����/�#U��������Nҭ�:˿�r��:����٠�;��8��6���ޘ��/n�*���}���I�J��5��^ӂ��&)^/=е�<}�Q���<g�s������W~J3ҿ��CE� F�	�|�!?�v���h��҂`�XT��	�ٍr���v����/�A�����+˔��هaD�C�fH��D�C{T��ٜ҆�S��Uf�|cU� Զ�]م�*"E�� [�����]c�]T��{+!��6 �c\2�#5^0+/���T� -^��f�3 � l�t��z6��9cǨ���aH�7�|2,3�~�e��O�qX��F�Jb68Q��|�5�̎lH�����^��?;�o���	����/t�"�(��.�#1��ͅ�ޯ�݅��k���p�����4`��KQ��-�n:�����Z��Q����V���@{)/����6���N����rK�/�(S�ŊQs!.�B�"���8�=��T�<�Zպr�S vL�X'�� $Ef7Ya�3���ѹP�A�.�h���z�ə4g�c���y���(3���q:����	:����K*�;��-L��2`�2�U�~6'�j�<k�+2؁ca�E@0,��:�Qv��J��뗝�Ȉ�	����&�~���S��\WA�b"&��f�Z6���?3g��o��f�5!����T�'��p���E�����v�]���f+�N�5{�����0�x�&v-��K�������F�o���[bH>VG��6n)�����;�X<t�2�������F!��d�;AC:���k���Ky��A�t�L��^Gϟ��|�M�m̭�4��j]�Gv��.�����v'MM����2"�`ưkhw���#B�kF/�qh7M����P>���(��1��eq�{�,�mzi��<jU�'w	��g�ejj��K3�z�+7=�0�rEX�c���p��u3d禯�k��f'Sؠ�s4
�ز[����[�V\���M�k����.r�_PY����?4���u��)X�{m-?�Ы�__J��'�ve�*"���%�4�t&u�O霢�:�T��9��?H[�u��7�2�2�$����7#s�1&����_q��x1~�Bԯ���yt��I�V�9 'K���cE�#V^z�pХ���=O��Ri�Ayv͗��g3�<�I�M�q��8����S���Q�6n�˭������s83`�z��C����d:��V$6̉	�swV�EV��"�F���^�~�Ըv2t�������.|bS�T�1|S^X��n�Х���хo+q��|���~xGl���۳Q�:�dp6˄�K�$r�� ��{6��-n���l<~>[:��Ә~����+�	=��\� �2�����4�ګ)F[�n
^��`ˍS���K��j���G�������C0i�Dƒy1C�P��#�t��+V�ڌ5x^�ݟo.���c(�DD�# �g��-�4�T��r��,�eF�/�n���g��A� 9��3���^U��:�p�MŦ�H����cl�)ݚ2^Y�w;V�s�{�8�a�����K[��MA_������40¾-<���;���'�sx{hԆ����]]h]N�8��/6���6o��S�F^Z��Y��0 �29��#Y%�*�MeH���#��N�y��JN�� �^���v���a3z��I�ɖ���ed�&��Hw|dd��|�m]�T��&ޥ��=������ϳ�7����Ұ�Oq"����>Z�7�K��RO�ߑ'���썪�ǐ�R}&�9x�)Z�	,���-cos���T7��������[	�H���*��M8�e�9E�5M#V��W��˒�s�?�����S�����N'=ک����8�,c%0�B��r�x�9��(��s�`��5�q��Iu�� p��>"��_�5/���;�&Q���%���a�U��,�O2�\�h}�v�kNu㥥��I�͈���b�3�V��P9QW'��P�
{�(쒔�>|�:����c��<��q�*Q6�3J�-nw(�[x��M�v�L��#K�6�w�w�������3PG�6��qIg��1_%���{�m�W��Y(py���,�}	H�ß9c4�$���X0�20�ݝ\��ŷy�9]�؜�̀�i�M�\�|_?�i�gY���%���qΩ��X���]���p�ЙB�<��P�ImL6EYv��3ߴ����"9�#�1�T���8%���2ݺ~>ˉ1S�f�I�3f{Q~�g�t�F��b�[P����C ���|�ka'p�R�y|���J�S
��,�t�X�nO�]	X�����J zG���Y�9�V�Y)��yt}$���B6`į*Dޛ5�c���,��V(�wx�Z ޾���r��ssc�vU*֦O`-O`]F��������3��xԆc��(��a8��e�	`�!�`�}���ƪ�w�� R:&x>�}�dp�oʊ$U�a�A_x�w���0���J3`_��$���%���댦���;	�� '�E�=蠽g��gp�'�feyK7�x��G!c�S(�d�n��z*,��4Q����EQq�˰H\�J��K>����,<��>ʷ�Ernk�ة/�&� W1w����<��usc�_��$�J�D�k����I��aR�a�׮&q�4+�\"���F�AB$��A<h. ����
�euvz}V�RT;a�L�r�,�8 /^^㢙C�I�R0%A�-��u��z��SCo� ��QI�B/�t��:��L�x�$U�ߦ
���E�7����f�M�>@�����g�d�+�ۅx�R��gV�Q�ۋ�\ԣ�G�:�.���;7��-��8}�Xt�)��$�ky������W�/���4�@��K����>��3{I���S�� Sc�SQ����F6���B�YmK����������C����!�O;�'�#t@}��0ni<m=f�f�@�B|�9���'�gz�*�-s&�q%��FQZ� /NM�?��,� ���b�[���[�@s��Ν	K���V��o�uIXTP��o �qu���N���.� �q�q����e��bwiEߊ��x��\l�u�tG*�l�}zy���_o/�ډ�媦2U� ���o���ݎ�-t3l<U����e�礱?U�ˠy�b��*�v�jq��%�HV�х<�^�1���[n��Ɖ��P߁��#�Vo��ޖ�
o����-��'ص��fsU��$�]��{�4�m)��WN~l�̋*�p�NK�8��H�
�5�ɀ�-{H�CE��֧��'>�`V�ٿ��a5��{�;�zP7���CMS8e���UZ�i�E���uA�|]����*~˸�"�A/����H��dЪr�U��K�^Ko�c���h|������G�3�����K����Рz���F�\��>���n"��`*��}N�|��*�
����|�%`���9D��Qe�F'����l�oV1�Ӣ�+R�G��e7�Q�]8}�9ߙ��0�x����nu�1�>�
��Jgs��g��<UV@՟Մz'�B�+2�+~��z�0�RQ��7١��U�&;{?QP��F0.�ժDM�[^��G9,�]�ll�k�(�ԥs!�+]XШ�����x���!���!     IEND�B`�PK   �K�X���DA  ~$     jsons/user_defined.json�ko�6��J�ϡ��%߆d����݀!H�l�9�+�+�b�}G��4��H^�h� �u�K�yyx�5[�/Bv�����)B,�Pd��_�Y�u'p�sG�k�^��N������޵�^����?����k���U�T7�py���M��j���yh����Y�v�|��>fQz0v(F��J��(G�X
!�b�7ga�r��v��8t�;�#�$"�C\;�L�yG"#�}��>�}�k[�M�.���΅�d�ɢ�ΫXg'_�j}wV.s{Z�!�ΩT��㩋�K{��\KIŶ�m��U�y��΋�US�2ķ��^��ޕs8"YΙ���smh��\�T�ۺ����U���ͭ�����>�/@t+ ��@7%�*ФPP�����
l@Av
b�O*��U d��H*�ލA�P�I9���1�
*��脙�I�W��i_ǄLxZMR�(`�6�<K�$r{��i�Nb�T���`���Q=f�Ik����k:F"�5��NBv��c$�`�=d�$Ĕ�H�M�������#�F��a{'���E�m���2i��ݝ�� i�� �����}��Ai�inuP����ݧ[4�4�7��zli�o��[DMN����L��	�}��A^Hӈ�>�� K�i�i�qu��DӐ�>����1gC�OJXt6��|��IgC�OJ��@�>���쓥YgC�OJ�Yv6��� K�Άh���ai����vfi���6�,<~�M)����>����4��;?H"M;��.�ćL� ֯7���m��Kلd�ES/B�*�ZPW@Zn;p�Uۢ�ݢj�Hv�n�]�b�I��˫l[����|�N�Ń~[�X.K7ǚ�y�Q�=�Q�m��֯�Mh�Q��8�����ն�c��h���qL9�>dDQ`�J��
Lt�*T���������k�mW��������6l��i���˙�R�;����My��.��٧���j�*���xtuAZ�Jn�Ҧ�f����1�\sd��0�
�ٱ7K�ZAZJ�Y���!���D�I��1�JQFQ�D�(*�^����2"5%aw�@��+u@���^�N�}M��i�sm��P��B���<-�]�~6�L��:�&'�?�5��r3K�}�A�a�3#�s����Մ�C�D��Qɞk�����<jm�B���]�oߧ��_������7ig�/��cg`#�^������Y�h�����h߶f��[�Vu��M].l�g\W��c��J����]�DLG�Xk$\�b��r'H\P�e �66 -����2j�taw�4d%"�T)��ID.�:�I`$����5,*�g���}/yl_l�y�a����7�!�B�I
SJ���s.q2F{�Kf1��+D�����7�꥓��g�R�%,����IE��`L�a�~�$�߹�6.8�ÎHY.P� _�(9���c݀+���(�A�i 7�N�)]h^���~,7(���ဤl3�C�]2��\ǐB�_� ���H��AG$��HK[��̍u��ǰyC2�n�1+k�I6� �n��?�p'�w< ���u��G�Ga�
BYr�\��PK
   �K�XЪ^-�&  kv                  cirkitFile.jsonPK
   J�X�R�� $� /             '  images/179c08ce-6e18-4019-8002-932a24469ad1.pngPK
   J�X��� �@ /             U� images/3e1f5452-c6ea-49ae-85fb-ddf6f8b38dad.pngPK
   J�X'(�5W �@ /             � images/4737cce6-ef6b-4e79-82eb-dab57378d86e.pngPK
   J�Xh`Pҷ!  �!  /             Y7
 images/4b60cb4e-ac73-4aba-afdc-1cf5937e57a1.pngPK
   ��X|�K�?  :  /             ]Y
 images/7720185d-ee5e-407b-a613-fa89a316821e.pngPK
   ��X��@��  ֈ  /             �n
 images/a2085874-a866-43e2-ad0b-af370f9f341d.pngPK
   J�X��t��"  �"  /             J�
 images/b09c32a2-0684-44ec-93cb-6718b830271d.pngPK
   J�Xr�>�� � /             f images/b24f041f-17b3-48b1-9f28-cb1f31b050cc.pngPK
   J�XF��-$  ($  /             r� images/d88a5b0e-66b3-4edb-b452-47f46dd40326.pngPK
   J�X?��O�o  �o  /             � images/ffe61187-e64a-4024-8cee-95dd034d2257.pngPK
   �K�X���DA  ~$               &� jsons/user_defined.jsonPK      $  ��   